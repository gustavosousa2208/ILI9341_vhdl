--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.07
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Thu Dec 15 12:07:39 2022

library IEEE;
use IEEE.std_logic_1164.all;

entity sprites is
    port (
        dout: out std_logic_vector(1 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(14 downto 0)
    );
end sprites;

architecture Behavioral of sprites is

    signal lut_f_0: std_logic;
    signal lut_f_1: std_logic;
    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_dout: std_logic_vector(0 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout: std_logic_vector(1 downto 1);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout: std_logic_vector(1 downto 0);
    signal dff_q_0: std_logic;
    signal gw_gnd: std_logic;
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);

    -- component declaration
    component LUT2
        generic (
            INIT: in bit_vector := X"0"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic
        );
    end component;

    -- component declaration
    component LUT3
        generic (
            INIT: in bit_vector := X"00"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic
        );
    end component;

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    prom_inst_1_dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    prom_inst_2_dout(1 downto 0) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    lut_inst_0 : LUT2
        generic map (
            INIT => X"2"
        )
        port map (
            F => lut_f_0,
            I0 => ce,
            I1 => ad(14)
        );

    lut_inst_1 : LUT3
        generic map (
            INIT => X"20"
        )
        port map (
            F => lut_f_1,
            I0 => ce,
            I1 => ad(13),
            I2 => ad(14)
        );

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F0077FFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_01 => X"FF1FF7F77FFFF7FFF7EFF7EFFFEFFFFF3FF7F77FE007E007EFF7E007E007FF7F",
            INIT_RAM_02 => X"EFFFFF7FF7F77FFFF7FFF7EFF7EFFFEFFFFF7FF7F77FFFF7FFF7EFF7EFFFEFFF",
            INIT_RAM_03 => X"EFFFEFFFFF7FF7F77FFFF7FFF7EFF7EFFFEFFFFF7FF7F77FFFF7FFF7EFF7EFFF",
            INIT_RAM_04 => X"EFFFEFFFFFF7FF7FF7F77EE007E007E007E007E007FF7FF7F77EFFF7FFF7EFF7",
            INIT_RAM_05 => X"EFFFEFFFEFFFFFF7FF7FF7F77EEFF7EFFFEFFFEFFFFFF7FF7FF7F77EEFF7EFFF",
            INIT_RAM_06 => X"EFF7EFFFEFFFEFFFFFF7FF7FF7F77EEFF7EFFFEFFFEFFFFFF7FF7FF7F77EEFF7",
            INIT_RAM_07 => X"FF7EE007E007EFFFE007E007FC1FF0077EEFF7EFFFEFFFEFFFFFF7FF7FF7F77E",
            INIT_RAM_08 => X"FFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_09 => X"FFFFFFFFFF7FFFFFFDFFFBFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0A => X"F7EFF7EFF7EFFF7FFFFFFDFFFBFFE007E007E007E0077FFFFFFDFFFBFFFFFFFF",
            INIT_RAM_0B => X"F7FFF7EFF7EFF7EFFF7E0001FDF80007FFF7EFF7EFF7EFFF7FFFFFFDFFFBFFFF",
            INIT_RAM_0C => X"FBFFF7FFF7EFF7EFF7EFFF7FFEFFFDFBFFF7FFF7EFF7EFF7EFFF7FFEFFFDFBFF",
            INIT_RAM_0D => X"FFFDFBFFF7E007E007E007EFFF7FFEFFFDFBFFF7FFF7EFF7EFF7EFFF7FFEFFFD",
            INIT_RAM_0E => X"7FFEFFFDFBFFF7EFF7EFFFEFF7EFFF7FFEFFFDFBFFF7EFF7EFFFEFF7EFFF7FFE",
            INIT_RAM_0F => X"EFFF7EFEFFFDFBFBF7EFF7EFFFEFF7EFFF00FEFC01FBFBF7EFF7EFFFEFF7EFFF",
            INIT_RAM_10 => X"E007EFFF7EFEFFFDFBFBF7EFF7EFFFEFF7EFFF7EFEFFFDFBFBF7EFF7EFFFEFF7",
            INIT_RAM_11 => X"FFFFFFFFFFFF7EFEFFFDFBFBF7FFFFFFFFFFFFFFFF7EFEFFFDFBFBF7E007EFFF",
            INIT_RAM_12 => X"000FDFDFBFBF007E7EFEFFFDFBFBF7FFFFFFFFFFFFFFFF7EFEFFFDFBFBF7FFFF",
            INIT_RAM_13 => X"FBFFFFFFDFDFFFBFFF7E7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFE01FC03FBF0",
            INIT_RAM_14 => X"FDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFF",
            INIT_RAM_15 => X"FEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFF",
            INIT_RAM_16 => X"FE7EFEFDFDF8000000001FC000007F007EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7E",
            INIT_RAM_17 => X"FF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7F",
            INIT_RAM_18 => X"DFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFF",
            INIT_RAM_19 => X"FFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDF",
            INIT_RAM_1A => X"F7FFEFDFDFFFBF7FFE7E00FDFC0003F00FEFDFDF803F007E7FFEFDFDFFFFF7FF",
            INIT_RAM_1B => X"FFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFB",
            INIT_RAM_1C => X"FDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFF",
            INIT_RAM_1D => X"7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFF",
            INIT_RAM_1E => X"FFFE7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFE00000003F7F0001FC03FBF0000",
            INIT_RAM_1F => X"BFBFFFFE7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFFFDFFFFFFF7FFEFFFDFBFBF",
            INIT_RAM_20 => X"FFDFBFBFFFFE7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFFFDFFFFFFF7FFEFFFDF",
            INIT_RAM_21 => X"F00FC01FBF80007E7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFFFDFFFFFFF7FFEF",
            INIT_RAM_22 => X"FFF7FFEFFFDFFFBFFF7EFEFFFDFDFFFFF7FFEFFFDFFFBFFF7E7E00FDFC000007",
            INIT_RAM_23 => X"FDFFFFF7FFEFFFDFFFBFFF7EFEFFFDFDFFFFF7FFEFFFDFFFBFFF7EFEFFFDFDFF",
            INIT_RAM_24 => X"FFFDFDFFFFF7FFEFFFDFFFBFFF7EFEFFFDFDFFFFF7FFEFFFDFFFBFFF7EFEFFFD",
            INIT_RAM_25 => X"FF7EFEFFFDFBFFFFFFEFFFFFBFBFFFFFFEFFFDFDFFFFF00FEFC01FFFBF007EFE",
            INIT_RAM_26 => X"BFFFFE7EFEFFFDFBFFFFFFEFFFFFBFBFFFFF7EFEFFFDFBFFFFFFEFFFFFBFBFFF",
            INIT_RAM_27 => X"FFBFBFFFFF7EFEFFFDFBFFFFFFEFFFFFBFBFFFFF7EFEFFFDFBFFFFFFEFFFFFBF",
            INIT_RAM_28 => X"0000003F8000007EFEFFFDFBFFFFFFEFFFFFBFBFFFFF7EFEFFFDFBFFFFFFEFFF",
            INIT_RAM_29 => X"FFFFEFFFFFFFFFFFFE7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFE0001F8000000",
            INIT_RAM_2A => X"FBFFFFFFEFFFFFFFFFFFFE7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFFFFFFFBFF",
            INIT_RAM_2B => X"FFFFFBFFFFFFEFFFFFFFFFFFFE7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFFFFFF",
            INIT_RAM_2C => X"7E00000003FBF00FEFC0000000007E7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFF",
            INIT_RAM_2D => X"FFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE",
            INIT_RAM_2E => X"FFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFF",
            INIT_RAM_2F => X"DFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFF",
            INIT_RAM_30 => X"FFFFDFFFFFBFFFFE0000FC01F803F7F00FDFC0000000007FFFFDFFFFFBF7FFEF",
            INIT_RAM_31 => X"FFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7",
            INIT_RAM_32 => X"FDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFB",
            INIT_RAM_33 => X"FEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFF",
            INIT_RAM_34 => X"7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E00FE01FDFBF807FFE000003FBF007E7F",
            INIT_RAM_35 => X"BF7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F",
            INIT_RAM_36 => X"FFFFBF7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E7FFFFFFDFBFFF7FFEFDFFFFF",
            INIT_RAM_37 => X"0FDFC0003F7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E7FFFFFFDFBFFF7FFEFDF",
            INIT_RAM_38 => X"FFFFEFFFDFFFBFFF7E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFE0001FBFBF000",
            INIT_RAM_39 => X"FBFBFFFFEFFFDFFFBFFF7E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFFFDFFFBFB",
            INIT_RAM_3A => X"FDFFFBFBFFFFEFFFDFFFBFFF7E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFFFDFF",
            INIT_RAM_3B => X"7E00FC000000000FE01FDFBF80007E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFF",
            INIT_RAM_3C => X"FFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE",
            INIT_RAM_3D => X"BFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFF",
            INIT_RAM_3E => X"DFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFF",
            INIT_RAM_3F => X"F7EFFFDFBFFF7FFE7EFE00000003F7F00FDFDF800000007EFEFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F0077FFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_01 => X"FF1FF7F77FFFF7FFF7EFF7EFFFEFFFFF3FF7F77FE007E007EFF7E007E007FF7F",
            INIT_RAM_02 => X"EFFFFF7FF7F77FFFF7FFF7EFF7EFFFEFFFFF7FF7F77FFFF7FFF7EFF7EFFFEFFF",
            INIT_RAM_03 => X"EFFFEFFFFF7FF7F77FFFF7FFF7EFF7EFFFEFFFFF7FF7F77FFFF7FFF7EFF7EFFF",
            INIT_RAM_04 => X"EFFFEFFFFFF7FF7FF7F77EE007E007E007E007E007FF7FF7F77EFFF7FFF7EFF7",
            INIT_RAM_05 => X"EFFFEFFFEFFFFFF7FF7FF7F77EEFF7EFFFEFFFEFFFFFF7FF7FF7F77EEFF7EFFF",
            INIT_RAM_06 => X"EFF7EFFFEFFFEFFFFFF7FF7FF7F77EEFF7EFFFEFFFEFFFFFF7FF7FF7F77EEFF7",
            INIT_RAM_07 => X"FF7EE007E007EFFFE007E007FC1FF0077EEFF7EFFFEFFFEFFFFFF7FF7FF7F77E",
            INIT_RAM_08 => X"FFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_09 => X"FFFFFFFFFF7FFFFFFDFFFBFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0A => X"F7EFF7EFF7EFFF7FFFFFFDFFFBFFE007E007E007E0077FFFFFFDFFFBFFFFFFFF",
            INIT_RAM_0B => X"F7FFF7EFF7EFF7EFFF7E0001FDF80007FFF7EFF7EFF7EFFF7FFFFFFDFFFBFFFF",
            INIT_RAM_0C => X"FBFFF7FFF7EFF7EFF7EFFF7FFEFFFDFBFFF7FFF7EFF7EFF7EFFF7FFEFFFDFBFF",
            INIT_RAM_0D => X"FFFDFBFFF7E007E007E007EFFF7FFEFFFDFBFFF7FFF7EFF7EFF7EFFF7FFEFFFD",
            INIT_RAM_0E => X"7FFEFFFDFBFFF7EFF7EFFFEFF7EFFF7FFEFFFDFBFFF7EFF7EFFFEFF7EFFF7FFE",
            INIT_RAM_0F => X"EFFF7EFEFFFDFBFBF7EFF7EFFFEFF7EFFF00FEFC01FBFBF7EFF7EFFFEFF7EFFF",
            INIT_RAM_10 => X"E007EFFF7EFEFFFDFBFBF7EFF7EFFFEFF7EFFF7EFEFFFDFBFBF7EFF7EFFFEFF7",
            INIT_RAM_11 => X"FFFFFFFFFFFF7EFEFFFDFBFBF7FFFFFFFFFFFFFFFF7EFEFFFDFBFBF7E007EFFF",
            INIT_RAM_12 => X"000FDFDFBFBF007E7EFEFFFDFBFBF7FFFFFFFFFFFFFFFF7EFEFFFDFBFBF7FFFF",
            INIT_RAM_13 => X"FBFFFFFFDFDFFFBFFF7E7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFE01FC03FBF0",
            INIT_RAM_14 => X"FDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFF",
            INIT_RAM_15 => X"FEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFF",
            INIT_RAM_16 => X"FE7EFEFDFDF8000000001FC000007F007EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7E",
            INIT_RAM_17 => X"FF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7F",
            INIT_RAM_18 => X"DFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFF",
            INIT_RAM_19 => X"FFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDFDFFFFF7FFE7FFEFDFDFFFFF7FFFFDF",
            INIT_RAM_1A => X"F7FFEFDFDFFFBF7FFE7E00FDFC0003F00FEFDFDF803F007E7FFEFDFDFFFFF7FF",
            INIT_RAM_1B => X"FFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFB",
            INIT_RAM_1C => X"FDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFF",
            INIT_RAM_1D => X"7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFFFDFFFFFBF7FFEFDFDFFFBF7FFE7EFF",
            INIT_RAM_1E => X"FFFE7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFE00000003F7F0001FC03FBF0000",
            INIT_RAM_1F => X"BFBFFFFE7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFFFDFFFFFFF7FFEFFFDFBFBF",
            INIT_RAM_20 => X"FFDFBFBFFFFE7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFFFDFFFFFFF7FFEFFFDF",
            INIT_RAM_21 => X"F00FC01FBF80007E7EFFFDFFFFFFF7FFEFFFDFBFBFFFFE7EFFFDFFFFFFF7FFEF",
            INIT_RAM_22 => X"FFF7FFEFFFDFFFBFFF7EFEFFFDFDFFFFF7FFEFFFDFFFBFFF7E7E00FDFC000007",
            INIT_RAM_23 => X"FDFFFFF7FFEFFFDFFFBFFF7EFEFFFDFDFFFFF7FFEFFFDFFFBFFF7EFEFFFDFDFF",
            INIT_RAM_24 => X"FFFDFDFFFFF7FFEFFFDFFFBFFF7EFEFFFDFDFFFFF7FFEFFFDFFFBFFF7EFEFFFD",
            INIT_RAM_25 => X"FF7EFEFFFDFBFFFFFFEFFFFFBFBFFFFFFEFFFDFDFFFFF00FEFC01FFFBF007EFE",
            INIT_RAM_26 => X"BFFFFF7EFEFFFDFBFFFFFFEFFFFFBFBFFFFF7EFEFFFDFBFFFFFFEFFFFFBFBFFF",
            INIT_RAM_27 => X"FFBFBFFFFF7EFEFFFDFBFFFFFFEFFFFFBFBFFFFF7EFEFFFDFBFFFFFFEFFFFFBF",
            INIT_RAM_28 => X"0000003F8000007EFEFFFDFBFFFFFFEFFFFFBFBFFFFF7EFEFFFDFBFFFFFFEFFF",
            INIT_RAM_29 => X"FFFFEFFFFFFFFFFFFE7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFE0001F8000000",
            INIT_RAM_2A => X"FBFFFFFFEFFFFFFFFFFFFE7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFFFFFFFBFF",
            INIT_RAM_2B => X"FFFFFBFFFFFFEFFFFFFFFFFFFE7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFFFFFF",
            INIT_RAM_2C => X"7E00000003FBF00FEFC0000000007E7EFFFFFFFBFFFFFFEFFFFFFFFFFFFE7EFF",
            INIT_RAM_2D => X"FFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE",
            INIT_RAM_2E => X"FFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFF",
            INIT_RAM_2F => X"DFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFFFFFFFFFE7FFFFDFFFFFBF7FFEFDFFF",
            INIT_RAM_30 => X"FFFFDFFFFFBFFFFE0000FC01F803F7F00FDFC0000000007FFFFDFFFFFBF7FFEF",
            INIT_RAM_31 => X"FFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7",
            INIT_RAM_32 => X"FDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFB",
            INIT_RAM_33 => X"FEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFFFDFBFFF7FFFFDFFFFFBFFFFE7FFEFF",
            INIT_RAM_34 => X"7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E00FE01FDFBF807FFE000003FBF007E7F",
            INIT_RAM_35 => X"BF7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F",
            INIT_RAM_36 => X"FFFFBF7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E7FFFFFFDFBFFF7FFEFDFFFFF",
            INIT_RAM_37 => X"0FDFC0003F7F7E7FFFFFFDFBFFF7FFEFDFFFFFBF7F7E7FFFFFFDFBFFF7FFEFDF",
            INIT_RAM_38 => X"FFFFEFFFDFFFBFFF7E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFE0001FBFBF000",
            INIT_RAM_39 => X"FBFBFFFFEFFFDFFFBFFF7E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFFFDFFFBFB",
            INIT_RAM_3A => X"FDFFFBFBFFFFEFFFDFFFBFFF7E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFFFDFF",
            INIT_RAM_3B => X"7E00FC000000000FE01FDFBF80007E7EFFFDFFFBFBFFFFEFFFDFFFBFFF7E7EFF",
            INIT_RAM_3C => X"FFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE",
            INIT_RAM_3D => X"BFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFF",
            INIT_RAM_3E => X"DFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFF",
            INIT_RAM_3F => X"F7EFFFDFBFFF7FFE7EFE00000003F7F00FDFDF800000007EFEFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"FF3FFF3FFCFFFFFFF3FFCFFFFFFF3FFFFFFC3FFFFFFCFFFFFFF3FFFFFFCFFF3F",
            INIT_RAM_01 => X"FFCFFF3FFF3FFCFFFFFFF3FFCFFFFFFF3FFFFFFC3FFFFFFCFFFFFFF3FFFFFFCF",
            INIT_RAM_02 => X"FFFFFFCFFF3FFF3FFCFFFFFFF3FFCFFFFFFF3FFFFFFC3FFFFFFCFFFFFFF3FFFF",
            INIT_RAM_03 => X"FFF3FFFFFFCFFF3FFF3FFCFFFFFFF3FFCFFFFFFF3FFFFFFC3FFFFFFCFFFFFFF3",
            INIT_RAM_04 => X"FFFFFFF3FFFFFFCFFF3FFF3FFCFFFFFFF3FFCFFFFFFF3FFFFFFC3FFFFFFCFFFF",
            INIT_RAM_05 => X"FFFCFFFFFFF3FFFFFFCFFF3FFF3FFCFFFFFFF3FFCFFFFFFF3FFFFFFC3FFFFFFC",
            INIT_RAM_06 => X"3FFC0000FFF3FFF3FFCFFFCFFF3FFF3FFC00000003FFC0000FFF3FFF3FFC3FFF",
            INIT_RAM_07 => X"3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFFFFFFFCFFFFFFF3FFF3FFC",
            INIT_RAM_08 => X"3FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFFFFFFFCFFFFFFF3FFF",
            INIT_RAM_09 => X"FFFF3FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFFFFFFFCFFFFFFF",
            INIT_RAM_0A => X"CFFFFFFF3FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFFFFFFFCFFF",
            INIT_RAM_0B => X"FFFFCFFFFFFF3FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFFFFFFF",
            INIT_RAM_0C => X"FFFFFFFFCFFFFFFF3FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFFF",
            INIT_RAM_0D => X"00FFF3FFF0000FFFC0003FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFF",
            INIT_RAM_0E => X"FFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFC0003FFF00000000000000000",
            INIT_RAM_0F => X"FFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFFFFF3FFFFFFFFFFFFFFFF",
            INIT_RAM_10 => X"FFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFFFFF3FFFFFFFFFFFF",
            INIT_RAM_11 => X"FFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFFFFF3FFFFFFFF",
            INIT_RAM_12 => X"FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFFFFF3FFFF",
            INIT_RAM_13 => X"FFF3FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFFFFF3",
            INIT_RAM_14 => X"FFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFC3FFCFFFF",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000000000000000000003FFC"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ad(14),
            CLK => clk,
            CE => ce
        );

    mux_inst_2: MUX2
        port map (
            O => dout(0),
            I0 => prom_inst_0_dout(0),
            I1 => prom_inst_2_dout(0),
            S0 => dff_q_0
        );

    mux_inst_5: MUX2
        port map (
            O => dout(1),
            I0 => prom_inst_1_dout(1),
            I1 => prom_inst_2_dout(1),
            S0 => dff_q_0
        );

end Behavioral; --sprites
