--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.07
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Tue Dec 13 01:03:24 2022

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(17 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(14 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal lut_f_0: std_logic;
    signal lut_f_1: std_logic;
    signal lut_f_2: std_logic;
    signal lut_f_3: std_logic;
    signal lut_f_4: std_logic;
    signal lut_f_5: std_logic;
    signal lut_f_6: std_logic;
    signal lut_f_7: std_logic;
    signal lut_f_8: std_logic;
    signal lut_f_9: std_logic;
    signal lut_f_10: std_logic;
    signal lut_f_11: std_logic;
    signal lut_f_12: std_logic;
    signal lut_f_13: std_logic;
    signal lut_f_14: std_logic;
    signal lut_f_15: std_logic;
    signal lut_f_16: std_logic;
    signal lut_f_17: std_logic;
    signal lut_f_18: std_logic;
    signal lut_f_19: std_logic;
    signal promx9_inst_0_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_0_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_1_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_1_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_2_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_2_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_3_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_3_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_4_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_4_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_5_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_5_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_6_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_6_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_7_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_7_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_8_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_8_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_9_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_9_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_10_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_10_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_11_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_11_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_12_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_12_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_13_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_13_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_14_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_14_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_15_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_15_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_16_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_16_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_17_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_17_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_18_dout_w: std_logic_vector(17 downto 0);
    signal promx9_inst_18_dout: std_logic_vector(17 downto 0);
    signal dff_q_0: std_logic;
    signal dff_q_1: std_logic;
    signal dff_q_2: std_logic;
    signal dff_q_3: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_11: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_13: std_logic;
    signal mux_o_14: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_31: std_logic;
    signal mux_o_32: std_logic;
    signal mux_o_33: std_logic;
    signal mux_o_34: std_logic;
    signal mux_o_35: std_logic;
    signal mux_o_36: std_logic;
    signal mux_o_37: std_logic;
    signal mux_o_39: std_logic;
    signal mux_o_52: std_logic;
    signal mux_o_53: std_logic;
    signal mux_o_54: std_logic;
    signal mux_o_55: std_logic;
    signal mux_o_56: std_logic;
    signal mux_o_57: std_logic;
    signal mux_o_58: std_logic;
    signal mux_o_60: std_logic;
    signal mux_o_73: std_logic;
    signal mux_o_74: std_logic;
    signal mux_o_75: std_logic;
    signal mux_o_76: std_logic;
    signal mux_o_77: std_logic;
    signal mux_o_78: std_logic;
    signal mux_o_79: std_logic;
    signal mux_o_81: std_logic;
    signal mux_o_94: std_logic;
    signal mux_o_95: std_logic;
    signal mux_o_96: std_logic;
    signal mux_o_97: std_logic;
    signal mux_o_98: std_logic;
    signal mux_o_99: std_logic;
    signal mux_o_100: std_logic;
    signal mux_o_102: std_logic;
    signal mux_o_115: std_logic;
    signal mux_o_116: std_logic;
    signal mux_o_117: std_logic;
    signal mux_o_118: std_logic;
    signal mux_o_119: std_logic;
    signal mux_o_120: std_logic;
    signal mux_o_121: std_logic;
    signal mux_o_123: std_logic;
    signal mux_o_136: std_logic;
    signal mux_o_137: std_logic;
    signal mux_o_138: std_logic;
    signal mux_o_139: std_logic;
    signal mux_o_140: std_logic;
    signal mux_o_141: std_logic;
    signal mux_o_142: std_logic;
    signal mux_o_144: std_logic;
    signal mux_o_157: std_logic;
    signal mux_o_158: std_logic;
    signal mux_o_159: std_logic;
    signal mux_o_160: std_logic;
    signal mux_o_161: std_logic;
    signal mux_o_162: std_logic;
    signal mux_o_163: std_logic;
    signal mux_o_165: std_logic;
    signal mux_o_178: std_logic;
    signal mux_o_179: std_logic;
    signal mux_o_180: std_logic;
    signal mux_o_181: std_logic;
    signal mux_o_182: std_logic;
    signal mux_o_183: std_logic;
    signal mux_o_184: std_logic;
    signal mux_o_186: std_logic;
    signal mux_o_199: std_logic;
    signal mux_o_200: std_logic;
    signal mux_o_201: std_logic;
    signal mux_o_202: std_logic;
    signal mux_o_203: std_logic;
    signal mux_o_204: std_logic;
    signal mux_o_205: std_logic;
    signal mux_o_207: std_logic;
    signal mux_o_220: std_logic;
    signal mux_o_221: std_logic;
    signal mux_o_222: std_logic;
    signal mux_o_223: std_logic;
    signal mux_o_224: std_logic;
    signal mux_o_225: std_logic;
    signal mux_o_226: std_logic;
    signal mux_o_228: std_logic;
    signal mux_o_241: std_logic;
    signal mux_o_242: std_logic;
    signal mux_o_243: std_logic;
    signal mux_o_244: std_logic;
    signal mux_o_245: std_logic;
    signal mux_o_246: std_logic;
    signal mux_o_247: std_logic;
    signal mux_o_249: std_logic;
    signal mux_o_262: std_logic;
    signal mux_o_263: std_logic;
    signal mux_o_264: std_logic;
    signal mux_o_265: std_logic;
    signal mux_o_266: std_logic;
    signal mux_o_267: std_logic;
    signal mux_o_268: std_logic;
    signal mux_o_270: std_logic;
    signal mux_o_283: std_logic;
    signal mux_o_284: std_logic;
    signal mux_o_285: std_logic;
    signal mux_o_286: std_logic;
    signal mux_o_287: std_logic;
    signal mux_o_288: std_logic;
    signal mux_o_289: std_logic;
    signal mux_o_291: std_logic;
    signal mux_o_304: std_logic;
    signal mux_o_305: std_logic;
    signal mux_o_306: std_logic;
    signal mux_o_307: std_logic;
    signal mux_o_308: std_logic;
    signal mux_o_309: std_logic;
    signal mux_o_310: std_logic;
    signal mux_o_312: std_logic;
    signal mux_o_325: std_logic;
    signal mux_o_326: std_logic;
    signal mux_o_327: std_logic;
    signal mux_o_328: std_logic;
    signal mux_o_329: std_logic;
    signal mux_o_330: std_logic;
    signal mux_o_331: std_logic;
    signal mux_o_333: std_logic;
    signal mux_o_346: std_logic;
    signal mux_o_347: std_logic;
    signal mux_o_348: std_logic;
    signal mux_o_349: std_logic;
    signal mux_o_350: std_logic;
    signal mux_o_351: std_logic;
    signal mux_o_352: std_logic;
    signal mux_o_354: std_logic;
    signal mux_o_367: std_logic;
    signal mux_o_368: std_logic;
    signal mux_o_369: std_logic;
    signal mux_o_370: std_logic;
    signal mux_o_371: std_logic;
    signal mux_o_372: std_logic;
    signal mux_o_373: std_logic;
    signal mux_o_375: std_logic;
    signal gw_gnd: std_logic;
    signal promx9_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_0_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_1_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_2_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_3_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_4_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_4_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_5_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_5_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_6_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_6_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_7_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_7_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_8_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_8_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_9_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_9_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_10_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_10_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_11_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_11_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_12_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_12_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_13_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_13_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_14_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_14_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_15_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_15_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_16_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_16_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_17_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_17_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_18_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_18_DO_o: std_logic_vector(35 downto 0);

    -- component declaration
    component LUT4
        generic (
            INIT: in bit_vector := X"0000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic
        );
    end component;

    -- component declaration
    component LUT2
        generic (
            INIT: in bit_vector := X"0"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic
        );
    end component;

    -- component declaration
    component LUT5
        generic (
            INIT: in bit_vector := X"00000000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic;
            I4: in std_logic
        );
    end component;

    --component declaration
    component pROMX9
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(35 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_gnd <= '0';

    promx9_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_0_dout(8 downto 0) <= promx9_inst_0_DO_o(8 downto 0) ;
    promx9_inst_0_dout_w(26 downto 0) <= promx9_inst_0_DO_o(35 downto 9) ;
    promx9_inst_1_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_1_dout(8 downto 0) <= promx9_inst_1_DO_o(8 downto 0) ;
    promx9_inst_1_dout_w(26 downto 0) <= promx9_inst_1_DO_o(35 downto 9) ;
    promx9_inst_2_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_2_dout(8 downto 0) <= promx9_inst_2_DO_o(8 downto 0) ;
    promx9_inst_2_dout_w(26 downto 0) <= promx9_inst_2_DO_o(35 downto 9) ;
    promx9_inst_3_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_3_dout(8 downto 0) <= promx9_inst_3_DO_o(8 downto 0) ;
    promx9_inst_3_dout_w(26 downto 0) <= promx9_inst_3_DO_o(35 downto 9) ;
    promx9_inst_4_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_4_dout(8 downto 0) <= promx9_inst_4_DO_o(8 downto 0) ;
    promx9_inst_4_dout_w(26 downto 0) <= promx9_inst_4_DO_o(35 downto 9) ;
    promx9_inst_5_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_5_dout(8 downto 0) <= promx9_inst_5_DO_o(8 downto 0) ;
    promx9_inst_5_dout_w(26 downto 0) <= promx9_inst_5_DO_o(35 downto 9) ;
    promx9_inst_6_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_6_dout(8 downto 0) <= promx9_inst_6_DO_o(8 downto 0) ;
    promx9_inst_6_dout_w(26 downto 0) <= promx9_inst_6_DO_o(35 downto 9) ;
    promx9_inst_7_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_7_dout(8 downto 0) <= promx9_inst_7_DO_o(8 downto 0) ;
    promx9_inst_7_dout_w(26 downto 0) <= promx9_inst_7_DO_o(35 downto 9) ;
    promx9_inst_8_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_8_dout(17 downto 9) <= promx9_inst_8_DO_o(8 downto 0) ;
    promx9_inst_8_dout_w(26 downto 0) <= promx9_inst_8_DO_o(35 downto 9) ;
    promx9_inst_9_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_9_dout(17 downto 9) <= promx9_inst_9_DO_o(8 downto 0) ;
    promx9_inst_9_dout_w(26 downto 0) <= promx9_inst_9_DO_o(35 downto 9) ;
    promx9_inst_10_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_10_dout(17 downto 9) <= promx9_inst_10_DO_o(8 downto 0) ;
    promx9_inst_10_dout_w(26 downto 0) <= promx9_inst_10_DO_o(35 downto 9) ;
    promx9_inst_11_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_11_dout(17 downto 9) <= promx9_inst_11_DO_o(8 downto 0) ;
    promx9_inst_11_dout_w(26 downto 0) <= promx9_inst_11_DO_o(35 downto 9) ;
    promx9_inst_12_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_12_dout(17 downto 9) <= promx9_inst_12_DO_o(8 downto 0) ;
    promx9_inst_12_dout_w(26 downto 0) <= promx9_inst_12_DO_o(35 downto 9) ;
    promx9_inst_13_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_13_dout(17 downto 9) <= promx9_inst_13_DO_o(8 downto 0) ;
    promx9_inst_13_dout_w(26 downto 0) <= promx9_inst_13_DO_o(35 downto 9) ;
    promx9_inst_14_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_14_dout(17 downto 9) <= promx9_inst_14_DO_o(8 downto 0) ;
    promx9_inst_14_dout_w(26 downto 0) <= promx9_inst_14_DO_o(35 downto 9) ;
    promx9_inst_15_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_15_dout(17 downto 9) <= promx9_inst_15_DO_o(8 downto 0) ;
    promx9_inst_15_dout_w(26 downto 0) <= promx9_inst_15_DO_o(35 downto 9) ;
    promx9_inst_16_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_16_dout(8 downto 0) <= promx9_inst_16_DO_o(8 downto 0) ;
    promx9_inst_16_dout_w(26 downto 0) <= promx9_inst_16_DO_o(35 downto 9) ;
    promx9_inst_17_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_17_dout(17 downto 9) <= promx9_inst_17_DO_o(8 downto 0) ;
    promx9_inst_17_dout_w(26 downto 0) <= promx9_inst_17_DO_o(35 downto 9) ;
    promx9_inst_18_AD_i <= ad(9 downto 0) & gw_gnd & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_18_dout(17 downto 0) <= promx9_inst_18_DO_o(17 downto 0) ;
    promx9_inst_18_dout_w(17 downto 0) <= promx9_inst_18_DO_o(35 downto 18) ;
    lut_inst_0 : LUT4
        generic map (
            INIT => X"0001"
        )
        port map (
            F => lut_f_0,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_1 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_1,
            I0 => ce,
            I1 => lut_f_0
        );

    lut_inst_2 : LUT4
        generic map (
            INIT => X"0002"
        )
        port map (
            F => lut_f_2,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_3 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_3,
            I0 => ce,
            I1 => lut_f_2
        );

    lut_inst_4 : LUT4
        generic map (
            INIT => X"0004"
        )
        port map (
            F => lut_f_4,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_5 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_5,
            I0 => ce,
            I1 => lut_f_4
        );

    lut_inst_6 : LUT4
        generic map (
            INIT => X"0008"
        )
        port map (
            F => lut_f_6,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_7 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_7,
            I0 => ce,
            I1 => lut_f_6
        );

    lut_inst_8 : LUT4
        generic map (
            INIT => X"0010"
        )
        port map (
            F => lut_f_8,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_9 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_9,
            I0 => ce,
            I1 => lut_f_8
        );

    lut_inst_10 : LUT4
        generic map (
            INIT => X"0020"
        )
        port map (
            F => lut_f_10,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_11 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_11,
            I0 => ce,
            I1 => lut_f_10
        );

    lut_inst_12 : LUT4
        generic map (
            INIT => X"0040"
        )
        port map (
            F => lut_f_12,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_13 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_13,
            I0 => ce,
            I1 => lut_f_12
        );

    lut_inst_14 : LUT4
        generic map (
            INIT => X"0080"
        )
        port map (
            F => lut_f_14,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_15 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_15,
            I0 => ce,
            I1 => lut_f_14
        );

    lut_inst_16 : LUT4
        generic map (
            INIT => X"0100"
        )
        port map (
            F => lut_f_16,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_17 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_17,
            I0 => ce,
            I1 => lut_f_16
        );

    lut_inst_18 : LUT5
        generic map (
            INIT => X"00040000"
        )
        port map (
            F => lut_f_18,
            I0 => ad(10),
            I1 => ad(11),
            I2 => ad(12),
            I3 => ad(13),
            I4 => ad(14)
        );

    lut_inst_19 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_19,
            I0 => ce,
            I1 => lut_f_18
        );

    promx9_inst_0: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"1C0DFEDB6DB5D1E26FD62A4CDA450564260CE9670D133DA8DCF0B99DDF27BBEDF6FB7DBE",
            INIT_RAM_01 => X"5CBEA773B9DCEE773B9DCEE773B9DCEE773B9DCEE7B3B9DCEDF73B9DBE9F6B95CAE47078",
            INIT_RAM_02 => X"5C2E572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B97D3EDF4FB",
            INIT_RAM_03 => X"9DCF77DBEDF6FB7DBE1C0D870761B1D86C351ADCEE772B95CF69B4DA0D86C763B2E170B9",
            INIT_RAM_04 => X"9DBE972B93C0E070381C7DB6D7499AC05FAC54AA348DFAC84C198A885644AF0DA8DCF0B9",
            INIT_RAM_05 => X"3C1E0F0FA7D4EDF53B9DCEEF93B9DCEEF93B9DCEE773BBE4EE773BBE4EE7B3B9DCF6773D",
            INIT_RAM_06 => X"DA0D46C363B2E170B85C2E170B85C2E0F0783C1E0F0783C1E0F0785C9E172B93C1E17278",
            INIT_RAM_07 => X"87A604A2EDA8DCF0B99DCF67BBEDF6FB7DBE1C1E0F0783C1E06C36DA5CEE532995CAE7B4",
            INIT_RAM_08 => X"9DCEE7B3B9ECEE773B7DAE572B91C0E3EE37FBEDAE935380BAD8A812895C159E962B8709",
            INIT_RAM_09 => X"3C1E0F0783C1E0F0383C1E172FA9DCEE773BBE4EEF93B9DCEE773B9DCEE773B9DCEE773B",
            INIT_RAM_0A => X"DA5CEE532994CAE573DA6D06A361B1D8EC763C1D8EC763B1E070783B0E06C381C1E0F078",
            INIT_RAM_0B => X"91179AF1184D0A068806A63482DDAFD8F0B99DCF77DBEDF6FB7DBE3C1E0F0783C1E0EC36",
            INIT_RAM_0C => X"9DDF2773B9DCEE773B9DCEDF4FB7D3EDF4FA5C9E0F0381C6DBEDF6DB4D666B0D6CA8CDE3",
            INIT_RAM_0D => X"1B0D86E361B0E070383C1E0F0783C0E06E373C3E9F4FA9DCEEF93BBE4EEF93B9DCEE777C",
            INIT_RAM_0E => X"3C1E172B93C1E0F036DA6D264F0993C265B4DA6D368351B0D8EC383B1D8EC381B0D86C36",
            INIT_RAM_0F => X"99AC45D291358941980A43A0F0240A050288A4A6349ADDAFD8F0FB9DDF37DBEDF6FB7DBE",
            INIT_RAM_10 => X"BE5F2777C9DCEE773B9DCEDF4FA7D4EE76FB7DBE9F6FA5CBED72B91C1E3EFF7FBEDB6D74",
            INIT_RAM_11 => X"1B0D86C761B0D86C361B0D86C36FB0D86E361C0D870383C0DC6E787D4EEF93BBE4EEF97C",
            INIT_RAM_12 => X"9DDF37DBEDF6FB7DBE5CAE572B95CAE57276DA5CEE532994CA6573DA6DB68351B0D86C36",
            INIT_RAM_13 => X"FBFDFEFB5DACCE66B037AA2B296C923812C8C23050200001010385A4857496CBA6D4F0B9",
            INIT_RAM_14 => X"9DCEE773BBE5F2F97C9DCEE773B9DCEE76FA9DBE9F4FA5CBEDF4FA5CAE572785C9E0F038",
            INIT_RAM_15 => X"B96D368351A8D46C361A8D86BB41A8D46A35DB6DB6DB6DA6D369B4DB6D36DF6DB0D8F0FA",
            INIT_RAM_16 => X"84A6249ADDAFD86EB99DCF77DBEDF6FB7DBE5CAE572B95CAE4EC361AED2E532783C5E373",
            INIT_RAM_17 => X"3C0E071F71BFDFEFB499CCCE02EB519A41DCE60188040A26148040200000000000008184",
            INIT_RAM_18 => X"994C9E332DB2E5F53B9DDF2773B9DCEE773B9DCEE773B9DCEE76FA7D3E972FB5CAE572B9",
            INIT_RAM_19 => X"1ADC9E0F0371B960F0994CAE772B9ED369B4DA6D36973B9CCEE532B94CA653278BC1E2F0",
            INIT_RAM_1A => X"41000000000000010244261422DBA6D4F0FA9DDF27BBEDF6FB7DBE7D2E572FA5CAE57076",
            INIT_RAM_1B => X"5C9E172383C0E3EFF7FB6DB6D35BA4CD606F1305292C1C2304808140D098400203058281",
            INIT_RAM_1C => X"170B85DEC16EB35BACD6EB05F335CCEE777C9DDF2773B9DCEE773B7D3E9F4FA7D3E9F6B9",
            INIT_RAM_1D => X"5CAE5F4FA5CAE57076DA5C85A2D157B05C6F379C160B0783C560B0582C16070381BCDE6F",
            INIT_RAM_1E => X"2010204004120582812010000000000000C102A6143ADDAFD86EB99DCF77DBEDF6FB7DBE",
            INIT_RAM_1F => X"7DAE572B95CAE4F0381C7DFEFB6BA5C9E0F037EB14010C66150281611008000613050240",
            INIT_RAM_20 => X"168B45A2DD66B2D56AB54AA552994AA150A8540B76CFA9DCEE773B9DCEDF6FA7D3E9F6FA",
            INIT_RAM_21 => X"9DCF67BBEDF6FB7DBE7D3E9F4FA7D2E57076B95C85BACD55AAD5ACD60B45A2E170B85C2D",
            INIT_RAM_22 => X"61205020040B0902402010184406120502C200100000000000008202A61422DDAED4F0B9",
            INIT_RAM_23 => X"7DAE572FA5CAE572783C0E0F038FB6DB6BB4589BFD9E40A93B0B850310080002020502C2",
            INIT_RAM_24 => X"168B45A2E170B85C2E168B85BADD66B3596C955AA552954AA5512916FD9F4FA9DBE9F4FA",
            INIT_RAM_25 => X"02A6248B1BA6D46EB99DDF27BBEDF6FB7DBE7D3E9F4FA7D3E97076B95C8542D155AB59AC",
            INIT_RAM_26 => X"C2C0902400000102C281B090200204090440408018440811010302200008040201008082",
            INIT_RAM_27 => X"1BAE5F4FA5CAE572B95C1E0F0383C0E3EE38FBEDB6974782C1606FF65B04C4E411010302",
            INIT_RAM_28 => X"3B5C9E06E168B85C6E373C1E0F0783C1E0F0782C160B0381C05A2D168B759EAD65AAD870",
            INIT_RAM_29 => X"0000000404110105020346648B1BA6D46EB99DCF6F9BEDF6FB7DBEBE3EAF8FA7D3E97076",
            INIT_RAM_2A => X"D64ABC7942010102C281C0D024020001030240C0E06812040D8481411020440811010344",
            INIT_RAM_2B => X"993C5E0F0383C1E2783C0DCF0783C7DF6DB4DA6DB6BB5DA6D2E9B4DA5D2E733582C0DE2E",
            INIT_RAM_2C => X"7D3E9F53B7D3E970B81A8D6E572783C2E572B9ED369B4DA6D369B4BA5CF6974B94CAE532",
            INIT_RAM_2D => X"81A06044060A050344200000040410008081036704B3399ED46EB97DCF67BBEDF6FB7DBE",
            INIT_RAM_2E => X"B94CEE533782C0DFACD64A7C759A230902C281C09048200101844040B098944813070AC1",
            INIT_RAM_2F => X"1B0D8F0361B0D46A35FB0D46BB4DA7D8F0B91B6DB69B4B9ED2E772B9DCAE773B9DCEE773",
            INIT_RAM_30 => X"7D4F77DBEDF6FB7DBEBE3EA773B7D4EE76B83B1D8EC35DA6DBEDF71B0D86C761B1D86C78",
            INIT_RAM_31 => X"81312894481C0A0744A230A88816120582C2201008081000000082446735B33DAFD8F0B9",
            INIT_RAM_32 => X"B9DD36974BA5D2E974BA5CA6532582C05DACB52A3499C4420503036240D8481408020944",
            INIT_RAM_33 => X"3C1E0F0783C2E572785C1E172783C1E0F0B83B0D86C361B9E1F437DB6D2E77399DCEE973",
            INIT_RAM_34 => X"06C8563B5DAED46EB97DCEE7BBEDF6FB7DBE9DBEA777C7D3EA76FA5C2E0EC351B0E07038",
            INIT_RAM_35 => X"40C0E050260A0480826240F09036240A07856140F0AC28130984C240A088082001000082",
            INIT_RAM_36 => X"FBEDAE773B9DCEE573B95CEE97399DCAE97399CCDE132581BC5DAC952A2C59AC620502C1",
            INIT_RAM_37 => X"5C9E0F0783C0E070781C1E170785CAE572B95CAE4F0B93C1E172B95C2E4F0783C2E5F4B9",
            INIT_RAM_38 => X"413088000202090282CA5B163B599FD8F0B97DCF77DBEDF6FB7DBEBE3EAF8FABE3E9F4FA",
            INIT_RAM_39 => X"952A245DC4820589846130985448140E888181512054460C0E8984A15128903A240D82C1",
            INIT_RAM_3A => X"5CAE0F0783C3EDF4B91C6DB6933BA5D2E532B94CE677299DCA6732994C960B1379BFD92A",
            INIT_RAM_3B => X"9DBE9F4FABE3EAF8FA5C2E070781B8E0F0781C1E0F0785CAE570B95CAE172B95C9E172B9",
            INIT_RAM_3C => X"C2D120503C240E04C2814090240002040104CE2C66733DAFD8F0787D4F67BBEDF6FB7DBE",
            INIT_RAM_3D => X"993C560B0378BB596A5489AC5DC081010503A22050281C2019850381D1206C260D120785",
            INIT_RAM_3E => X"5CAE570B95C9E172B93C2E4F0785CBE9F4FA1C1E07037DB6DB697299DCA6733B94CE6532",
            INIT_RAM_3F => X"7D4F67BBEDF6FB7DBEBE5F2F8FABE3E9F4FA5CAE0EC783C0DCF0783C1E0F0785CAE572B8"
        )
        port map (
            DO => promx9_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => promx9_inst_0_AD_i
        );

    promx9_inst_1: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"40D1206C16101B0B84C2D1308C281C0A88C2A26108082202090448508BE6735DAED4F0B9",
            INIT_RAM_01 => X"DB5D2E93399CCA66F078AC1606F177B3592A5489A45DB48101028181611848181E1606C2",
            INIT_RAM_02 => X"3C1E0F0783C2E572B95CAE4F0B95C1E172B85CAE4F0785CCEDF4FA3C2E0F0383C0E3EDB4",
            INIT_RAM_03 => X"B62C66733DAED4F0B97DCEE7BBEDF6FB7DBE9DBEA76FABE3EAF8FA5C2E0F0383C0E0F038",
            INIT_RAM_04 => X"8140A0681818160702815130902810180D84C2C0C0D44813068902826150200411010488",
            INIT_RAM_05 => X"7D2E572785C9E07038FBFDB6DB4BA4CE6732992C5606F176B2D8E83369645DBC62050281",
            INIT_RAM_06 => X"5C2E0F0363C1E0F0783C1E0F0B93C1E172B85CAE572B95CAE172B95CAE4F0787D3EA76FA",
            INIT_RAM_07 => X"8140D020040901051917BCDE733DAED4F0FA7DCF67BBEDF6FB7DBEBE5F2F97CBE3EA76FA",
            INIT_RAM_08 => X"33692439A8490103444130A8902A26140B84A26130B02A20180D44623070B85812060503",
            INIT_RAM_09 => X"5CAE4F0B97DCEE76FA5CAE572FA5CAE572B93C0E3EC37DB6DAE933993C4DE6F176B254A8",
            INIT_RAM_0A => X"BE5F2F97C7D4EE76FA5C2E0F0783C1E0F0373C1E0F0783C1E172B95C2E4F0B95C9E172B9",
            INIT_RAM_0B => X"A240A06068130A07038140902824100209A5D6CCE66F3DAFD8F0B99DCEE7BBEDF6FB7DBE",
            INIT_RAM_0C => X"DA4CD6270D66B254E8136914159C24088082C2A060744620140B8502E130B44036130B85",
            INIT_RAM_0D => X"5CAE570B95C9E172B95CAE4F0787D3E9F4FA7DAE4F0B95CAE572B95CAE4F0381B8DFEFB5",
            INIT_RAM_0E => X"7DCEE7BBEDF6FB7DBE9DDF2777C9DDF276FA5C9E0EC783C1E0F0783C1E0F0B93C1E172B9",
            INIT_RAM_0F => X"C2E160606C2B128985C240A07858240A890360E12048160800902D17BCDE73399FD86EFA",
            INIT_RAM_10 => X"7D2E572781C0E071F6BA4CDE0B016EB254A8F25894119A220984814120A058481D120785",
            INIT_RAM_11 => X"3C1E0F0783C1E172B95C2E570B95CAE570B95CAE4F0B97D3E9F6FA5C9E172B95CAE572FA",
            INIT_RAM_12 => X"17BC9E533DAED4F0B97DDF27BBEDF6FB7DBEBE5F2F93B9DCEE76FA5C2E170783C1E0F037",
            INIT_RAM_13 => X"40A090303C240A0784A250A8985035130848C2C0E8805C2C0B0B448130A048260A06282F",
            INIT_RAM_14 => X"7D1E0F0B93C2E572B97D2E572B93C0E3EFF6DB5D1E26F16EB254A8F2489C01540A050240",
            INIT_RAM_15 => X"5CAE0F0783C1E0F0783C1E0F0783C1E172B95CAE4F0B85CAE572B95C9E172785CBE9F4B9",
            INIT_RAM_16 => X"81C120882814081BAD58AC56333DAFD86EB97DCF77DBEDF6FB7DBEBE4EE777C9DDF1F4FA",
            INIT_RAM_17 => X"F1C883A0D40A05024040A050481C2E118303A101B0A05035100A060340A0544C240A8944",
            INIT_RAM_18 => X"5CAE172B95CBE9F6B95C9E172B93C2E572B95CAE572B93C0DC6FF6DB5D264B1176B1D026",
            INIT_RAM_19 => X"9DCEE773B9DDF1F4FA5C2E4F0783C1E0F0783C1E0F0B95C9E172B85CAE172B95CAE570B9",
            INIT_RAM_1A => X"02C0B0984C2C0E0503C2205050282306236C58BCDE6F2DA8DCF0B97DCEEF9BEDF6FB7DBE",
            INIT_RAM_1B => X"DA6D664B016DAA5226D248BB80681511048140A050542A251204C26140E8806035100B85",
            INIT_RAM_1C => X"5CAE572B85C9E172B95CAE572B97D3E972785C9E0F0781C1E070B91C1E0F0381B0DC71F6",
            INIT_RAM_1D => X"7DCF67BBEDF6FB7DBE9DCEEF93B9DCEDF4FA5CAE4F0783C1E0F0783C2E4F0783C1E0F0B9",
            INIT_RAM_1E => X"61206898503513080602C0C0B44C25118282A22050302414082B6C58AC562F3DAED5F4FA",
            INIT_RAM_1F => X"3C0E06FF7DB0DC71B699CCD626FF66B15226B1486328140C0A048240B090584C230606C2",
            INIT_RAM_20 => X"3C1E172785C9E172B95CAE172B95C9E172B95CAE570B97D2E572B93C0E070381C0E07078",
            INIT_RAM_21 => X"17BC96333DA8DCF0FA9DCF67BBEDF6FB7DBE9DCEEF93B9DCEE76FA7D2E4F0783C2E4F078",
            INIT_RAM_22 => X"4140A0503C2C0A8944811000B840350B098502E130B03C2C0903028120502C14140AA56C",
            INIT_RAM_23 => X"1C0DC71F71BFDFEFF6FB7DBEC36DB7DB6DB5BA4CD6270D65A95026B1286A4812010104C2",
            INIT_RAM_24 => X"7D2E572783C1E0F0785C9E0F0783C2E0F0785CAE572B95CAE172B93C2E572FB5CBE97278",
            INIT_RAM_25 => X"81205028260A06236C58AC562F3DAED4F0FA7DCF6F9BEDF6FB7DBE9DBE9F53B7D4EDF4B9",
            INIT_RAM_26 => X"9117B18C18130800402020880C2C2512890281A068903036170805C26128903C2C0A0584",
            INIT_RAM_27 => X"3C2E572FA5CBE97278FB8DC6DF6FB0DC6DB6BA6DB6DB5DB7DBED74BA4CDE06FD64A95068",
            INIT_RAM_28 => X"7D3E9F73B7D3E9F4FA5CAE4F0783C2E5F4783C1E0F0783C1E170785CAE4F0B95C2E570B9",
            INIT_RAM_29 => X"0351288C2A240E040641205028161205112917BC9E4F2DA8DCF0FA7DCF67BBEDF6FB7DBE",
            INIT_RAM_2A => X"99CCD606FD65B15226916711144A230A064020102054240D130902C2D130985C2E128806",
            INIT_RAM_2B => X"3C2E570B95CAE172B95CAE572FB7D9E070381B8DBEDB6FB6DB69B4DA5CAE974DA7DB6D74",
            INIT_RAM_2C => X"9DCF6F9BEDF6FB7DBE7D3E9F4FA7D3E972B95CAE4F0B93C1E172783C2E4F0783C1E17278",
            INIT_RAM_2D => X"02E130985A240985854451182C18140A0544612060440412040D2917AC562F3DAED4F0B9",
            INIT_RAM_2E => X"99CCE6572DB6DB6BB4BA4CD606F16DB1D1E49126309038140E0682202060544C2C0A8903",
            INIT_RAM_2F => X"5C9E0F0783C1E0F0785C1E0F0B95CAE570B95CAE572FB5C9E07038FBEDB6BB5DA5D26733",
            INIT_RAM_30 => X"B60BD62F3DAED4F0B99DDF27BBEDF6FB7DBE5CAE572B95CAE572B95C2E4F0785C9E0F078",
            INIT_RAM_31 => X"8161504400351308C1A2015118581A0585854440E05448130A08C14120502812020B08A9",
            INIT_RAM_32 => X"DB6DB6D74BA5CAE732995CA67B4DB7DB6D74BA4CDE26F176B152265003584C14090184C1",
            INIT_RAM_33 => X"5C9E0F0783C1E172783C1E0F0783C1E0F0785C9E170B95C9E172B95CAE572FB5C8E071F7",
            INIT_RAM_34 => X"C2411050240C12049FB62C562F3DAFD8F0B97DCF6F9BEDF6FB7DBE7D3E972FA5CBE972FA",
            INIT_RAM_35 => X"2F42502406130903448140B088140E1708C1C25121385C240B0A062440905044140A0902",
            INIT_RAM_36 => X"5CAE5F6FA5C8E0F1F7FB6D36974995CAE53258CCEE9F6FBEDB6DB6BA4CD626F175A95026",
            INIT_RAM_37 => X"5CAE572B95CAE572B95C9E172785C9E172785C9E0F0783C1E0F0783C1E172B95C1E172B9",
            INIT_RAM_38 => X"8140A0984818191088032200B04A2122881554AC562B1DAFD86EFA9DCF67BBEDF6FB7DBE",
            INIT_RAM_39 => X"99BC56070D64A84D228CD1104400010185038120689444140A8806818151185C2C0E8984",
            INIT_RAM_3A => X"3C1E0F0B95CAE570B95CBE9F4B95C9E06FF6DB6DAE9B499CCA64B0994CFEC37FB7DB6B74",
            INIT_RAM_3B => X"9DCF6F9BEDF6FB7DBE7D3E972B95CAE572FA3C2E572B93C1E0F0783C1E0F0783C1E0F078",
            INIT_RAM_3C => X"C26100D850340B0AC2A26130903C65241B8C06E31100660A22881012EB45EB199FD86EB9",
            INIT_RAM_3D => X"BA7DBEC38FB5D36974992C0DE2ED63A3C8E006A0A050240B0502820340E0405A23040D84",
            INIT_RAM_3E => X"3C1E0F0783C1E0F0783C1E0F0783C2E172B97D2E5F4B93C0E3EDF7DB6D2E733994CA66F1",
            INIT_RAM_3F => X"0EDB05EF299ED4F0FA9DCF67BBEDF6FB7DBE5CAE572B97D2E572B95C9E172B95CAE57278"
        )
        port map (
            DO => promx9_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => promx9_inst_1_AD_i
        );

    promx9_inst_2: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"410170805036130805C26130B84C230A08C144527180D0865228900AC442109028180B09",
            INIT_RAM_01 => X"FBEDAE73399CCA6774FB7DBEDF6FB6DAE933580BB5BAC741A2C5DC81A090502811020481",
            INIT_RAM_02 => X"5CAE572B95CAE4F0B93C1E0F0783C0E0F0783C1E0F0785CAE172B97D3E972B91C0E06DB6",
            INIT_RAM_03 => X"0AE51304E484081A064C5B05EB19AED572FA9DCF6F9BEDF6FB7DBE7D2E5F4B95CAE572FA",
            INIT_RAM_04 => X"4100080C1614098584C240E89028481A880502D100D84036151184848341A90272623319",
            INIT_RAM_05 => X"7D3ED72781C0DBEFB6DB4D6E933B9ED369F61BFDBEDF6DB5D266F1378B7592A336954098",
            INIT_RAM_06 => X"5CAE572B95CAE572B95C9E1F4B93C1E0F0783C1E0F0783C1E0F0783C1E0F0785C9E172B9",
            INIT_RAM_07 => X"A4C262352A8855419CCE155AE150AA41214DC62A75A2FDAED572FB9DCF67BBEDF6FB7DBE",
            INIT_RAM_08 => X"D65AA52A812E913E05202098584408020744812200C88C2221118424613080684A200A0D",
            INIT_RAM_09 => X"3C1E172783C2E572785CAE572381C7DB6DB5DA5D2E974BA6D76C371B7DFEDF7BA3C45C2E",
            INIT_RAM_0A => X"9DCF77DBEDF6FB7DBE5CAE572B95CAE572B95CAE5F4785CAE4F0783C1E0F0783C1E0F078",
            INIT_RAM_0B => X"036130A8823446124E87830AA554B05541215007931596B8542A9088AA6D82F999E1F4FB",
            INIT_RAM_0C => X"1BFDB6D74991BC5DACD64A4CC26D23823344000010281815130B44A20140A064401A1206",
            INIT_RAM_0D => X"3C1E0F0783C1E0F0783C1E0F0B95CAE4F0B95CAE4F038FBFDB6D74BA6D6E974DB7D86E36",
            INIT_RAM_0E => X"4C262D9ADDA8DD72FB9DDF2F9BEDF6FB7DBE5CAE572B95CAE4F0B95CAE572785C9E0F078",
            INIT_RAM_0F => X"A26100B85032211109034261307A493AA5526B955AF92CD46749A4F1870385EEE056B39C",
            INIT_RAM_10 => X"DB6DA67B5BA7D86E38FB4CDE270F66B2D52A542A44C26913802A4000000808240E100A05",
            INIT_RAM_11 => X"3C1E0F0783C1E0F0783C1E0F0783C1E172785CBE8F0785C9E0F0B93C1E0F037FBFDBEDB6",
            INIT_RAM_12 => X"7066941DB2F281C01D5087551ACDA8DDF4FA9DCF67BBEDF6FB7DBE5CAE572785C9E0F078",
            INIT_RAM_13 => X"408000081813070B03811188C05E2A208D0902C249D09C90321FDCCD4623194CD0784DA4",
            INIT_RAM_14 => X"DB0DCF078FBFDBED35BA6D76BB6FB7DBED74780B85DAC953A1D0A9330984C25B12822282",
            INIT_RAM_15 => X"3C1E0F0785C9E0F0785C9E172785C9E0F0783C1E0F0783C2E4F0783C0DBEDB4B92C2666F",
            INIT_RAM_16 => X"EE771AE5C4F48B485E0E07A405E0F28244A1502815070DA8DD72FB9DCF67BBEDF6FB7DBE",
            INIT_RAM_17 => X"1309BC9A4912801A4000101040040C0F0A064440D91494441D1006A4C1F280DE9549B159",
            INIT_RAM_18 => X"587B358E873AA04520AF2A358B0995D36D74BA5D2E974BA4CD622DD64A14CA833298CC26",
            INIT_RAM_19 => X"7DCF67BBEDF6FB7DBE5CAE4F0783C2E4F0783C1E0F0783C1E0F0783C1E0F0783C7DA66F0",
            INIT_RAM_1A => X"87834191087E49AE1E707692D185078CBDDA90489405ED109A45210EE92522FDA8DD72FA",
            INIT_RAM_1B => X"3209849E4F189049E3F1F9349627017A88000040D0205232228806C64248C06C562A9311",
            INIT_RAM_1C => X"3C1E0F078FB0BE64B0F61BAD4A8120923C9D8B66741A2114ABD82E583C5E2F1588BA54A8",
            INIT_RAM_1D => X"1299950B1DA8DD72B99DDF2F9BEDF6FB7DBE3C1E0F0B93C1E0F0783C1E0F0783C1E0F078",
            INIT_RAM_1E => X"C52389D0927033288EA943EA2148804E321E7066B25182F6883C5C9007AC52270486441D",
            INIT_RAM_1F => X"732A3586E175A84C669178EC320905864161B0E8A44E07077102000040B0A0583C1D1107",
            INIT_RAM_20 => X"3C1E0F0783C1E0F0783C1E0F078DAAC45CB0956AAC3A2D137F3399AA96B32DD2D57A4120",
            INIT_RAM_21 => X"900793DDC4C3804CA854CAAD974DA8DCF0FA9DCF77DBEDF6FB7DBE3C1E0F0783C1E0F078",
            INIT_RAM_22 => X"40A08810306E281B070613B15492754921940A25AA359C9050BC1E70278AAD80F1783C1C",
            INIT_RAM_23 => X"AAD54B5D629555BA956EE82BD694EC38259109299CF204F070381E6F9793C5EEE2600000",
            INIT_RAM_24 => X"3C1E0F0783C1E0F0783C1E0F0783C1E0F0373C1E0F078BA1C05A2F780B43529541993BD6",
            INIT_RAM_25 => X"6F871B118D1278B8DF2F079412250AA04CE8542A15333DA8DCF0FB9DCF6F9BEDF6FB7DBE",
            INIT_RAM_26 => X"CD566B21C0A138800060A058384C2222130784E289D0F87A3921514B750AA14884612C1C",
            INIT_RAM_27 => X"992A15066176913B55AAA5732528963B9D55292552B558F2943512AAE461CA65478F359A",
            INIT_RAM_28 => X"9DCF77DBEDF6FB7DBE3C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078DB2C3582E",
            INIT_RAM_29 => X"2AE69B01CA8A392D590E072B3DAB0F73C6A0ED992C5A4744A44C665419AD933DA9E0F0FB",
            INIT_RAM_2A => X"D62A23CA654690381C70565B19ACA5489000409028985028140C0683E2A0E0C88E291D92",
            INIT_RAM_2B => X"3C1E0F078FB3C65226333C7D826177933399AAE8333128914A15CEC7644A599124A741A0",
            INIT_RAM_2C => X"94CA85B33DA9E172FB9DDF27BBEDF6FB7DBE3C1E0F0783C1E0F0383C1E0F0783C0E0F078",
            INIT_RAM_2D => X"27443140C87A5B2414C964BB8D88804FB9DA91170389E2E27B4520F189345A5948984D2A",
            INIT_RAM_2E => X"4AA54A49DCCD579C07D0198CD6AD62A1CEE7335884DE4ACA4318C144222938C0370D918A",
            INIT_RAM_2F => X"3C1E070783C1E0F0783C1E0F078FB2C553E4F26A96066D62A3329DCCF9332D8EB03E15C7",
            INIT_RAM_30 => X"1268A4466D64A9536A533A153B5FB0DD72FA9ECF77DBEDF6FB7DBE3C1E0F0783C1E0F078",
            INIT_RAM_31 => X"2AE53155247139908EC94391D92A966AB214A90712D9288442A2D82F073349EACC83C9E3",
            INIT_RAM_32 => X"704A5B11EC89481F55D2230948C2930E0280C3683C624530915024952A2556A54382B352",
            INIT_RAM_33 => X"3C1E0F0783C1E070783C1E0F0783C0DCF0783C1E0F0783C5D1E1E45378F58A8D62A341A0",
            INIT_RAM_34 => X"0A564B89E6FC834520B0873C7ACB65AA53DC884635BB5DA8DD72FB9DDF27BBEDF6FB7DBE",
            INIT_RAM_35 => X"944AA54E8954A14DE44F17334D7A9752A214C543DB19206773B559AC871B0140A04CAAD8",
            INIT_RAM_36 => X"543805D2A95689C199D1382D2A8C894B1CDDD612909462914B83C1E051A2D918F171C120",
            INIT_RAM_37 => X"9DCF67BBEDF6FB7DBE3C1E0F0783C1E06E783C1E070783C0DCF0373C1E0F0783C0DEE928",
            INIT_RAM_38 => X"EE156B39A4B3602855A8973B69EB0C83C9202F792552A954A65120ED17B5933FB0DD72FA",
            INIT_RAM_39 => X"62E011580012564161944A5D0A694AA250E712793B9DCEE25829DB09A5AA5920A66B3559",
            INIT_RAM_3A => X"3C1E070783C1E2662E94688DDAC33585C1209517B549D4AA321C9DB4E3B8E8C466661D91",
            INIT_RAM_3B => X"950B85F331B8DCF0FA9DCF77DBEDF6FB7DBE1C1E0F0781B9E0F0783C0DCF0373C0DCF037",
            INIT_RAM_3C => X"4F383B9D48835F25182A84C38D8EA0512D92C966BB59AB0C8240DFD13A2D96A955AA5466",
            INIT_RAM_3D => X"3314894DD872584DA0C8E2509810117344A673A9A54A6D56A8CCA612790385C2E37C3855",
            INIT_RAM_3E => X"3C1E0F0783C0DCF0783C1E0F0783C1E06EB037AA0CDAC54099C1A254898CDDC4EE45CEA8",
            INIT_RAM_3F => X"124AB59ACD66B05C2D176B05F741B8DCF0FA9DCF77DBEDF6FB7DBE3C0DCF0783C1E0F078"
        )
        port map (
            DO => promx9_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_5,
            RESET => reset,
            AD => promx9_inst_2_AD_i
        );

    promx9_inst_3: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"D169349E3CD76B441E0E283C99A70051B19AED35F3455C9155AF182AE6B341C4F47B44DF",
            INIT_RAM_01 => X"172C3C8E04AF71A0E0F22558B994EF7151E4132578286C8890CCE794EABD5AAD539C4864",
            INIT_RAM_02 => X"1B8E0F0371B8DC6E371B8DC6E371B8DC6E371B8DC6E783C0DC6F33D2CAA452A344A93D2A",
            INIT_RAM_03 => X"2AE69BEDF6FC81BFE3B14AAD42E171BCDE2DF66B1E533FB1E172FA9EDF27BBEDF6FB7DBE",
            INIT_RAM_04 => X"F629A51AA9499A40DF739984DE32E25745E3B12A3489E0F079C19AED64A205587051AF9A",
            INIT_RAM_05 => X"379BF4AE054EB359AC954AB58D86EC80CD61D666723994E9984DE433584A495B0998CCE8",
            INIT_RAM_06 => X"9ECF77DBEDF6FB7DBE1BFD86E371B8DC6E37FB0DC6E371B8DC6FF6FB0DFEDF63C3E97238",
            INIT_RAM_07 => X"2E04F2520A8853359A8C0513C1C2E47A3C22334AB582E170B85BACD66B0E1B5FB0DD72FB",
            INIT_RAM_08 => X"33098449ED2299516AF639E5066F22A044A6946AB49A20E4392CDF903A3C8269007AC21E",
            INIT_RAM_09 => X"FB7DBEDF63C2E57237DB2C7581D504ABD9229499B589E6C753C866D6361B0E06C693592A",
            INIT_RAM_0A => X"952996333DA8DD72FB9DCF77DBEDF6FB7DBEFB7DBEDF6FB7D86FF6FB7DB6BF6DB7DBEDF6",
            INIT_RAM_0B => X"532A23C24D2199C05E0F64BB813EA4622DDA09E6A305CED0724120950B85C7037AA241A2",
            INIT_RAM_0C => X"D6585C0260E29A54261319B44A6542994CA6D56A94CE794299CEA6534A048964723AC2E8",
            INIT_RAM_0D => X"FB7DB6BF6FB6D7EDB5FB6D7EC373C3E9F678DACD6D9AC134AB59A5547924466CCA55B122",
            INIT_RAM_0E => X"740B4DEB0172A0AA1AEA15561B5FB1E172FB9DCF77DBEDF6FB7DBEFB7DBEDF6FB7DB6BF6",
            INIT_RAM_0F => X"B0873300A87170CCE8D63A048E0124A1CEE78C07241DC4B2793C1447172B214ED27A40DF",
            INIT_RAM_10 => X"D60924024EE773B8E094F9150264F0995026332A244A81329B5466B56AAD4E89539CCD28",
            INIT_RAM_11 => X"FB7D86FF6FB7D86FF6FB7DBEDF6FB7DBEDF6FB7DBEC785CBE972781BCCC5FACF26B244A0",
            INIT_RAM_12 => X"A8B5DB0D76C172409EB50BBD82D379BB596A386B0E1331B8DD72FB9DDF27BBEDF6FB7DBE",
            INIT_RAM_13 => X"D60B85D2A94383B813C884AB28E4B381D1AC16CA23D16112A358A8D1071C05C6FC5A1C13",
            INIT_RAM_14 => X"DB4CCE16CD62A2D86F54C8B3320700913DA4917904DE4F248950A8B52A05CA8956B16129",
            INIT_RAM_15 => X"9ECF77DBEDF6FB7DBE1B8DC6E371B8DC6E371BFD86FF61BFD86FF61B8DC6EB97DBE97238",
            INIT_RAM_16 => X"33198BCD70E068285CCC383559ACD1543920376B05CB1586B14C22126B163B5FB0DD72FB",
            INIT_RAM_17 => X"1309A552AD67B3546E170BAD56A2E25A200A09D47B9A20E2A2542E94CA03599D17AA552A",
            INIT_RAM_18 => X"1B8DCF0FA7D3E8F038DACCC5F6C0F0B95266176AAC320F22753CA8D25855266954A950A8",
            INIT_RAM_19 => X"C0871E5B5DA9E172FA9DDF37DBEDF6FB7DBE3C1E0F0783C1E06E781B8DC6E371B8DC6E37",
            INIT_RAM_1A => X"950682452324A7596A5309839A2ACD8744D7D125B3118D1564385C546B0DEB0385AA3C8D",
            INIT_RAM_1B => X"D61984CA8332A2552A744AA53AC54DABD9ACB52C05D2AB0E491B10475484D2AD60B7D82D",
            INIT_RAM_1C => X"3C0DCF0783C1E0F0781B9E172FB9DAE46FB69ACCD616A132875BAC914AB4A66F2199C066",
            INIT_RAM_1D => X"583C05C6F376B04998C8A61E7B5DA8DD72FB9DCF77DBEDF6FB7DBE3C1E0F0783C1E0F037",
            INIT_RAM_1E => X"4F39C5BECF60B45BAC5468A1D5EB50B45D6AB52A244E0D23803DDAACF6AB21C6F972B264",
            INIT_RAM_1F => X"B60984C2633690CD2A583A04CA8136B358E8F63A3596AD60BB596AF66B3596ACC443A9DC",
            INIT_RAM_20 => X"3C1E06E783C1E06E783C1E0F0783C1E0F0781B9E1F4FA7D2E7EFB6BA4CCDD6AD6CAA5529",
            INIT_RAM_21 => X"ACC8335DA2E27A31DB741BF596A176B05DECB50B5E5B5DA8DD72FB9DCF77DBEDF6FB7DBE",
            INIT_RAM_22 => X"D60BAD56A4F23BB92AD66AB592994EB05CE85376A2C24D60BBD9ACF64AB58A833099C05C",
            INIT_RAM_23 => X"BA2C5E2F0380BCD1AC54A804C26956944D6AD6EB1D1A4744AA532A5489BD8A8B53A359AC",
            INIT_RAM_24 => X"9DCF77DBEDF6FB7DBE3C0DCF0371B8DC6E371BFD86FF61B8DC6E371B9E172B93C7DFEFB6",
            INIT_RAM_25 => X"944A6D5A4D299A41DC9027A40DF4F37C3920133C0DE66D60B7582DD62A267B5FB0DDF4FA",
            INIT_RAM_26 => X"956B1D0A9742A45D2AD65AB592A4B0313DAC171B8DCA67329A546ED6544B520B56B05C2E",
            INIT_RAM_27 => X"FB1E172381C0DF6DB699CCE66F358AC6D868D607540A1334A953AC956B34B2A54CA951AC",
            INIT_RAM_28 => X"176B267B5DA8DD72FA9EDF27BBEDF6FB7DBEFB8D86E36FB7D86DF6FB7DBEDF6FB7DBEC35",
            INIT_RAM_29 => X"120722C24B56B3596A734A1D1ACB51993DDC0E768B86690278B99A132A6D5AC954A85C2E",
            INIT_RAM_2A => X"952A1532AD63A1D0A695099D129B54AB59AC170BA55292AC58482E173C0DDEA3229744E7",
            INIT_RAM_2B => X"DB6D769B5DAED36DB5DB2E47038DB6DB6D74BA6D26AF3999C35A26D22C358A9334A9D12A",
            INIT_RAM_2C => X"705A85D29B5790CC2ED66B267331B8DCF0FA9DCF77DBEDF6FB7DBEFB6DBEDB6DA6DB6BB4",
            INIT_RAM_2D => X"171B961AC52D7844E611478B824944A0DC6ED1093D4B0F669039D20E37C381C6C669BE9E",
            INIT_RAM_2E => X"4C56758E8336B3592A132A2D56AD66B151A4746B2552AF66B2542E170BB58E7EE27651EC",
            INIT_RAM_2F => X"BA5D2E97499DD2E933BA5D2677499DD2E933DA9E0F1F71BFDF6BB6FB6D76D3358EB655A4",
            INIT_RAM_30 => X"6C178399A11662B3DAB0A7A55AC950922C4E6C2A1E7B51B8DD72FB9DDF37DBEDF6FB7DBE",
            INIT_RAM_31 => X"D60B85C242E4A2553237FB3D8B073276BC22122765264746ABD56AB5088C9EAB52A24024",
            INIT_RAM_32 => X"FB6DB6B3317DB0D015886292DA4955A9D1AC546B1536AD67B254A8544A950E8D6199516A",
            INIT_RAM_33 => X"9DCF77DBEDF6FB7DBE99CCE673399CCE653399CCE673399CCE6772DB0E06FB6FBFDBEDF7",
            INIT_RAM_34 => X"73B9FD52853193C7200A688AB160D66B31181127A45AC9519B44D02AC61E3B5DA8DD72FB",
            INIT_RAM_35 => X"54EB151299527B496A16EB14D162AD49A0E0171B8DC2E7368340A51145A3D1E5408BD52A",
            INIT_RAM_36 => X"FB0DFEDF6DB7DBEFF7FB6D666B1956942B110A05329A4334AA55AC543A2C56AD6FB253AC",
            INIT_RAM_37 => X"4AA626BB5DA8DD72FB9DCF77DBEDF6FB7DBE99DD2673399CCE6532994CE673299CCE6774",
            INIT_RAM_38 => X"1106834229458AD5AC73891CE22534A94C1C1276A1C0A8F170389EB0B824466B55B255E3",
            INIT_RAM_39 => X"956B2D4A9546B150E8B55A84CA96FC614DECD60991AC1A6D3719424327B582E1508B411E",
            INIT_RAM_3A => X"99CCE653399CCE67B4FBFDB6DB6DB0E071F7DB4D667B0342A1AF188825BC762545B2452A",
            INIT_RAM_3B => X"D10904C26744AB592A5319A6774FB1E1F4FB9DCF77DBEDF6FB7DBEBA5D2E97499CCE6733",
            INIT_RAM_3C => X"A93052B283247A3C5A4EC5B4064947A85DAA950B445A0941984561C9170124E2AC613D59",
            INIT_RAM_3D => X"4B48231E43358950A9F62A6536AB609B48A95499952A8B0873D82ED661688C88704B22D7",
            INIT_RAM_3E => X"BA5D2E933B95CAE533B94CEE97299DD2E9B61BED36933DB0DFEFB6DB4CDE7AD13671AF0F",
            INIT_RAM_3F => X"1164B44140A259BF20F209245E45469255AC955AA67331B9E172FB9DCF77DBEDF6FB7DBE"
        )
        port map (
            DO => promx9_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_7,
            RESET => reset,
            AD => promx9_inst_3_AD_i
        );

    promx9_inst_4: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"4F715900DD84B904108813A851E53088355E0D1693A22533A05C2E954A848A5F509B441C",
            INIT_RAM_01 => X"9ACCC5E2FD2A812C14270784C66135AAD4A8137B2536A332A15026912A150662E4605B2A",
            INIT_RAM_02 => X"9ECF77DBEDF6FB7DBEB95CAE53399CCE673299CCAE53399DCAE9F6FB6D369B41C0DC6FB6",
            INIT_RAM_03 => X"375A9CFEA9429A401CC958735D22766839204F48344A6F1998486694098E1B5FB1E0F0FB",
            INIT_RAM_04 => X"952A6D9292E19A55AC441008C000000001044654510D0D5294B422AF1904520116ABD9EC",
            INIT_RAM_05 => X"1BED2E8371B8DFEDB69ACCCE16C91077B85547463345EEE58B48A8D26B35AA8D65AA53AC",
            INIT_RAM_06 => X"F209963331B9E1F4FB9ECF77DBEDF6FB7DBEB94CAE572995CA6572994CA6532995CAE9F6",
            INIT_RAM_07 => X"AAB984464900B45B6A94FB0CD28D50913CA68C668481CED565AF91CC275C1E3F1F8FC626",
            INIT_RAM_08 => X"F1AA2D52A950995068D2EB153AC5358551AC231008C000000001044154719CC33587AD1E",
            INIT_RAM_09 => X"994C9E332994CAE9F6DB6DB6A785C9E36B35998BED868CE27BC992A8C422C142E278481C",
            INIT_RAM_0A => X"EE48048E7131984DE4B0E92D9331B9E1F4FB9ECF77DBEDF6FB7DBE99BC5E33278CCA64F1",
            INIT_RAM_0B => X"825441AC812192BD160D27444DF326B0DC6E176B3D5EA7399B55DA8C154AAD709A3BA4D7",
            INIT_RAM_0C => X"50E9131612A95693206BA9A44E8500784C66134A45C2DD699B552A409031400000000084",
            INIT_RAM_0D => X"994CA653278CC9E332994CA6532995CAE9B61BED070B93C7DA66F317EB55226D2565219C",
            INIT_RAM_0E => X"ACB7E41590902A920C09F6F44A894893C8263379267331B9E1F4FB9EDF37DBEDF6FB7DBE",
            INIT_RAM_0F => X"608009D0F15210014DE925A08C8D139E1D55D008A3C220E0BB58B0371BBD8F05429AC29E",
            INIT_RAM_10 => X"9489A45228C99BB89691283B89EA8C59C11088A83B9DCD17703C1E1358A542DD67B3D82D",
            INIT_RAM_11 => X"9EDF37DBEDF6FB7DBE993C66532994CA64F1993C5E332995CA66361C0DDF4FB1C4CD616C",
            INIT_RAM_12 => X"331B8DE2ED67A8489E4F76A3198EA04C180A47462C26694CA5D1A51348951331B9E172FB",
            INIT_RAM_13 => X"CD5654362B65A9D16A06615831154C842916E9220008E53682AA22113984422C54CA55EC",
            INIT_RAM_14 => X"5C9E1F6FBFBAC45AE8F24803DA26BF71B1490A238AA2653079AFA2EE466A5CC0F278AAE0",
            INIT_RAM_15 => X"12793D9B51B9E172FB9ECF77DBEDF6FB7DBE994CA6532995CA657278DCA6532B95CAE837",
            INIT_RAM_16 => X"32680B5988B0B755AC372C3D82E174A8CDE34F072401CB0C8B240AE945BC6A894CA84C24",
            INIT_RAM_17 => X"0A024ABA28C565C0E82A857281CACEB05B2994F1401044813A2290240038ADFD514BAC22",
            INIT_RAM_18 => X"994CAE572BA5CB68375CAE676B9FB3C2D4669027A3151A895429226BD484920ACB81D0E7",
            INIT_RAM_19 => X"88438B824F2199CEA873F9355B61B9E1F4FB9EDF37DBEDF6FB7DBE993C6E532993C66532",
            INIT_RAM_1A => X"46204AB2915169BAE70D2291B20A88B5CEDFF60B9606FD65B1516211663B4DF2E278B8D7",
            INIT_RAM_1B => X"A487345DB7428244A86FF308C13C923A32E8B136220D06C17AD42ED50918302002110884",
            INIT_RAM_1C => X"994CAE4F1994CA6532995CAE572B95CB6A785CBEA76FA1B9C25426906682998E9239910E",
            INIT_RAM_1D => X"91171BF205037E41200A07331611339CCCA69419A55351BAE572FB9ECF77DBEDF6FB7DBE",
            INIT_RAM_1E => X"580BB4455E2B11040000256BD5EAF579CC5AC8C4B171ED16B2C529580B85C2E377B0CC66",
            INIT_RAM_1F => X"6F9733198471542992C964AB264D609A33ACB5382D424902A3B9A4370B75826F24A5506F",
            INIT_RAM_20 => X"9ECF77DBEDF6FB7DBEB93C6E532994C9E372994CAE572B96D368787D3EA76FA1BAC25226",
            INIT_RAM_21 => X"B50B7D9AC168BAD4A81219345A2D178DBE1E880722C1E134AAD529954A85DB51B9E1F4FB",
            INIT_RAM_22 => X"94EB6542F586B05CF0583C45C2EF256798C4E602A1D128975B9C47E71684495D13C3B62D",
            INIT_RAM_23 => X"5CBEE76FB1BBC75866F1A7BB718C93211C24D2793C9DC4C323340C6BBA0BD9287566A4F0",
            INIT_RAM_24 => X"B64AA55741B9E1F53BBE5F37DBEDF6FB7DBE994CA653278DCA6572784CAE532B95CAE878",
            INIT_RAM_25 => X"2D189CCA5780BB5572171BF582ED67B05AE85309048241278E41DACA442A3DA123A2552A",
            INIT_RAM_26 => X"8A19B4A261241E2D20EDEB04D6CB50985DECD62C1E2F017EB0B999EA0280DCC0A51A8DCE",
            INIT_RAM_27 => X"994CA6572B95CB68385CCEE76FB1C4CFD929F1A8231594AE492D8B8866A319A9107633E4",
            INIT_RAM_28 => X"4B170ABDAD13A1D1AC952A45BB51B8DDF4FB9EEFB7DBEDF6FB7DBE994CAE4F1994C9E372",
            INIT_RAM_29 => X"2D2751B9146A2A1D552D579CDEA996B3586E54EB358A6746B05DAC3309048241258A41DC",
            INIT_RAM_2A => X"4F66AA213ACA79C15254467B9ACD287A20952918B44E7177B04D28D54A04CA9D62C35424",
            INIT_RAM_2B => X"994CA6532B93C66532994CAE572B95CAE8377D4EE773B5CDD0E1AD3358BB6D7C92582951",
            INIT_RAM_2C => X"7409049E4F1C8BB759CD769BFA2132A2D52A94DAAD9331B8DDF4FBBE4F77DBEDF6FB7DBE",
            INIT_RAM_2D => X"947AAC4A6D57AB59AA94FB1CC5AC8A38130E29148C42D581B8DCB0B519A55E373DA85B6A",
            INIT_RAM_2E => X"9499BC7186BA3B160C09C834551A9071CF20A9567449EF1B9D204E0E68034E6175A8D0E7",
            INIT_RAM_2F => X"9EEFB7DBEDF6FB7DBE785CA64F0B94CA6572993C66532B95CB69F65CBEE773B5CFD9E22F",
            INIT_RAM_30 => X"D6299C1A273DA85BAC7389849E4F1C883855CA35F48A8743A2D4A812F9151331B9E172FB",
            INIT_RAM_31 => X"8819241982D6894DE313091CFA2122994BAA16CA1CC5A0543B230E8771722E7170B85D6A",
            INIT_RAM_32 => X"3C3EE773B7D8DEE6F1D6CA84BDC0A2591C14A8D27A8D770381900CACC6220D71137C1549",
            INIT_RAM_33 => X"542A15133DA9E1F4FBBE4F77DBEDF6FB7DBE994C9E132B93C5E132994CA6532B95CA67B5",
            INIT_RAM_34 => X"8711880D0331C3492A950993DA2944A759ACB54A5CEE712D883A964F68AC4A894CAAD4E8",
            INIT_RAM_35 => X"09E2A2110A4E4B878AE93050C0A2906A3C223208B446452B9D4DAAB54A5CD5EAA9491991",
            INIT_RAM_36 => X"784CA64F1995CAE574FB3E9F53B7D1E36D74386B759A4ACF4B17948B04C2949C907A4414",
            INIT_RAM_37 => X"EDE88CCA6744A9D12954CA65333FB1E1F4FB9EEFB7DBEDF6FB7DBE994CA64F0994CA6532",
            INIT_RAM_38 => X"94988C55E2D554B41A4AE1000864A9904C24F2383B422125A85DAC94AA0CC25F1B83B61C",
            INIT_RAM_39 => X"2746345D294652C50F8C5269286C56288C4609B20150E09168348A094792C5C32274C8A5",
            INIT_RAM_3A => X"783C1E0F0783C1E0F0783C264F0994CA6572DB2E5F4FA7D3EBEFB599BC75A25EE25B248E",
            INIT_RAM_3B => X"74097C65E2F5652C0C6F891D0E8954A654A8F21A359B5DA8DDF53BBE6FB7DBEDF6FB7DBE",
            INIT_RAM_3C => X"0F170C8E6D0088446473680B55BEB16B325A05306844060A57B4D8CCB613A64B55ABD9AC",
            INIT_RAM_3D => X"BA6D4E16CEE5651C960E285C1EC3358950E054589AEA02F6B2D425531562CE66F991BF1E",
            INIT_RAM_3E => X"9EEFB7DBEDF6FB7DBE783C1E0F0783C1E0F0783C1E132B94CA6533DA9E1F73B9DBE8F038",
            INIT_RAM_3F => X"4443834E6537A85A2D54790BC982AF6D3D2090090CCE8B55AA52A83469359B5DA9E1F53B"
        )
        port map (
            DO => promx9_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_9,
            RESET => reset,
            AD => promx9_inst_4_AD_i
        );

    promx9_inst_5: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"8714A2C2273AA2D522B519242665478CCC6411192BDD6EB554B5CE686178A86C2A089C15",
            INIT_RAM_01 => X"DA8DDF4FA7DBE972781BFDB6A2D1285739DC0F6903BAC344A84CA1B55A8CD62CD4463086",
            INIT_RAM_02 => X"541A359B51B8DDF53BBE4F77DBEDF6FB7DBE583C1E0B0782C160B0782C160B0994CA6733",
            INIT_RAM_03 => X"2971702C140A0881C564255BB1E940B85BAC5437FB79C2AF6FC66612093C6A83319A52E8",
            INIT_RAM_04 => X"336B2441206254B9E3332A04B2994CA4CD2A941994C26702A255AA7389045D6EB168B516",
            INIT_RAM_05 => X"582C160B0784CA653399FD9F4FA7D4EDF6B93C1E36CB0137505CA013771C159D10944D2A",
            INIT_RAM_06 => X"532984C24F1AA550A9544935B351B8DD733D9EEFB7DBEDF6FB7DBE782C160F0582C160B0",
            INIT_RAM_07 => X"335864095C8C592A95887150C88A1259B1DA46C5B4128D61B8DFACF24813194ED973C824",
            INIT_RAM_08 => X"EA7321C5EC92A241590EE2A2D1ED169359ACD60B4E16CF64A6D826949A2556A547B1CCE7",
            INIT_RAM_09 => X"582C160B0582C160B0582C1E0F0784CA673399ED4F0B97DBEDF6FA5C9E3ED3317BA3B952",
            INIT_RAM_0A => X"91773B855B0F8C4866331984DE4706904AA8344845BB51B8DD733B9EDF37DBEDF6FB7DBE",
            INIT_RAM_0B => X"B55CDD09E3269345A02D5561C0AC8E3A1D91E2A2317914EE8B45E42E171CDAAF60B85C26",
            INIT_RAM_0C => X"5C9E3ED74D6876239AA89551D922E35F24D787E481BC3D20944AA8547AB592A950B85D6A",
            INIT_RAM_0D => X"9EEFB7DBEDF6FB7DBE582C160B0582C160B0582C160B0583C6653399CD46EFA7D3EDF73B",
            INIT_RAM_0E => X"13278CC2ED60B952A191071C120D178FC666330904D22505643BA512E7255B51B9E1F53B",
            INIT_RAM_0F => X"06A61C122955A85C2F785ABC8DFEE651A0C8435090C4E46A2A1C8DA482B32A6952A550A8",
            INIT_RAM_10 => X"99CD7ECFA7DBEDF73B7D2E46F74D6876B2146BA7AC29E0E2782910F187034554ED442A4E",
            INIT_RAM_11 => X"0EC675BB53C1E1F53B9EEFB7DBEDF6FB7DBE582C160B0782C160F0582C160B0784CA6733",
            INIT_RAM_12 => X"D04AB582E37EB2D5AC95092502E377B150A0916693C24127914C2613792C5DC4FC652098",
            INIT_RAM_13 => X"1378C4920AC9541952A8E33482ED67B05DE44C2210440005369286A4E451546C4D54345A",
            INIT_RAM_14 => X"582C160B0783C6653399CD76CB99DBE9F6FB7D2E46F35B67703D20134A04D61535864120",
            INIT_RAM_15 => X"D15883B19A965212100AA6252373C3E9F73B9EEFB7DBEDF6FB7DBE583C1E0F0783C1E0F0",
            INIT_RAM_16 => X"F2189BB5545228B422948B8E02E580BB59ACB54AB582ED648942A0CD071BFE4F209849E4",
            INIT_RAM_17 => X"4F790CC26F62A04D6253199C1225048029DC6FE9653AC950B64584C2A2213094100204D8",
            INIT_RAM_18 => X"994CA6532994CA64F0582C1E0B0583C66533BA4D76A787DBED72FA7D2E46EF10ED66B3E4",
            INIT_RAM_19 => X"F24824026120904DA24F7722314080400C8844042D9B51BAE5F73D9EEFB7DBEDF6FB7DBE",
            INIT_RAM_1A => X"4FA67188E47534008E1129BAC9D2D43AAA95D1198DF2A582C05FEC168B45DAD3417941A4",
            INIT_RAM_1B => X"3C1E26B2A4B6481898134A84DAC542A242A91319A55E4D24894226D24A758E8541578A0C",
            INIT_RAM_1C => X"9EEFB7DBEDF6FB7DBE995CAE572B95CE6572783C1E0F0784CA673399DD36BF67DBECF078",
            INIT_RAM_1D => X"581BC5BAC54692C4A89529B44261209AC5627035D2006C2C1C1B0702C5255B51BBE9F73D",
            INIT_RAM_1E => X"B52A3496A136130B490000000820695511092E6B0A51EAF277AC0A2E66B58E8580B961AD",
            INIT_RAM_1F => X"99ED76BB63C3E972371BAC6C59C6C05244A1D66B1516A94BA151E454E9748A0B17913EA8",
            INIT_RAM_20 => X"27466D9B51BAE5F53B9EEFB7DBEDF6FB7DBEB95CAE772B9DCAE532994C9E0B078CCA6733",
            INIT_RAM_21 => X"8B48354E8176B560B0378BAD8A81309950A8742A150A81378EC25E505481B8403321118A",
            INIT_RAM_22 => X"D62A349A4914AB58A8F2483C8E80AD0A9200000000000412412040CC398B41A2E6883516",
            INIT_RAM_23 => X"B94CA64F0784CA6733BA6D36BB61BAE5723878EB03959EE098DD6C131A150A8131A1D0A8",
            INIT_RAM_24 => X"AC8500C46446289D9287C66D9741BBEA773D9EEFB7DBEDF6FB7DBEB9DCF6973B9ED2E773",
            INIT_RAM_25 => X"0E4A6AA5A110894B1E0E39DD12A581C1E06FD66B2D4A954099D12A54BA254A95438345DC",
            INIT_RAM_26 => X"0F2A1512A954AAD5A5911984C263419B58264F3A153A4272041200420000082426292040",
            INIT_RAM_27 => X"DA6D369B4DA6D36972B94C9E132994CE6733BA5D36BB6FB9E17278D6D88299C136B1432A",
            INIT_RAM_28 => X"953A152665448A441CE9238120A4684C2751A8C645B333C3E9F73DBE6FB7DBEDF6FB7DBE",
            INIT_RAM_29 => X"9278C00820343C8C86F22952B552D190C8E7900B85C66582C45C2EF65AAD5AC13198CCA9",
            INIT_RAM_2A => X"CE462442E168BA54A8B52A358A9954A84C25D6692452A54E97C762F2092D4E8E6207180D",
            INIT_RAM_2B => X"9EEFB7DBEDF6FB7DBEDA6D369B4DA6D369B4B9DCA6532994CA6733BA5D369B6FB8E06EB1",
            INIT_RAM_2C => X"D56B0CCA95489950A9544A44C2613488B81C0A648190EA8F482613870745F331BBE9F73D",
            INIT_RAM_2D => X"54198CD290F6169B0E875340C0DA8854808D13483301A11190C8A6C60B9E322170BB5928",
            INIT_RAM_2E => X"BA5D36BF6FB7DEE85E6B898DE2E582A04D2AD1790CDECD209AD522332A140663309BC826",
            INIT_RAM_2F => X"C94885F351BBE9F73DBE6FB7DBEDF6FB7DBE1AED06BB41A8D769B4B9DCA6532994CE6774",
            INIT_RAM_30 => X"CD0BA65A4D61BA50A8956B151E412E904DA4D2E934A2513488399A47238120A8804C2613",
            INIT_RAM_31 => X"952A13EA912E90CCE854AA6D52A9011903140AB5C2751A9615A1208F068341A4AF92552A",
            INIT_RAM_32 => X"DA5CAE532994CA6774BA6DB6DF6FBCCE42D7F60B953ACD64A8CC26B0C8049ACD60955226",
            INIT_RAM_33 => X"4B4622C55097491B0FA8F9163351BAE6773DDF6FB7DBEDF6FB7DBE3B0D86A351A8D46A35",
            INIT_RAM_34 => X"4AE80B4A60D08A536AD51BD622ED56B2D5EC132A44C261377142A1D24884D22D238230D8",
            INIT_RAM_35 => X"B09993DACF679150A9542A34AA8D219B5826134A8CC2654549A192821200C48E2F51602E",
            INIT_RAM_36 => X"1B0D86C363B0D46BB4B9DCEE532995CE6BB5DAEDBEDF61C280BC2ED60BB59ACD609B4529",
            INIT_RAM_37 => X"50282C5A490769AE1C4F76DAE9687748269509C89E7351BAE6777C9EEFB7DBEDF6FB7DBE",
            INIT_RAM_38 => X"332843C24D61B9CE5AAF06B412812296522DF62C1606ED64A05D6AD2095412450C66B25E",
            INIT_RAM_39 => X"131BD61ACD60B8CD201227B49AD955A8CCA91309950E854AA5532A742A6552A543813B22",
            INIT_RAM_3A => X"DF6FB7DBEDF6FB7DBE3C1D8EC763B1D8EC35DA5CEE532B95CAE9B4DAED86DB40E8B85D2A",
            INIT_RAM_3B => X"B548820980F54B2922913813CE0CD76A41206F8733095090492A95E9669E174FB2E6773D",
            INIT_RAM_3C => X"5409952A8B1649AFE4950BD606F37EB3449DF248045291219BC8A8379B960B0F66B255AC",
            INIT_RAM_3D => X"DB0DF6C68F63A160A8171B85DAC540B9506690682D92A37BA1526633097C8A9331A3592A",
            INIT_RAM_3E => X"09E71E535FB2E5F73DDF6FB7DBEDF6FB7DBE3C1D8F0763B1D8EC35DA5CEE57299DCAE9B5",
            INIT_RAM_3F => X"F57B05C2D955AB58E8B1672A415C9633299A50091BE1C6FE8B45A290772B3168B45A2C12"
        )
        port map (
            DO => promx9_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_11,
            RESET => reset,
            AD => promx9_inst_5_AD_i
        );

    promx9_inst_6: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"951A358E8134AA556C94CAA55E48C442B224D66B1602EF64AB41A01247AD2A8D068A51A2",
            INIT_RAM_01 => X"1ADCEE572B9DD369F6FBDCFD82E3719B58A8955B0DE26540BBC8A8D008B5A2D174AB5826",
            INIT_RAM_02 => X"EE66B35988B45A2D160956563331BBE9F73DDF6FB7DBEDF6FB7DBE5CAE172B93C1D8EC35",
            INIT_RAM_03 => X"122994B61CC88A3DA2915AA5529174A8CD215048B2911C662AA5184F37E40DFD109345A2",
            INIT_RAM_04 => X"6C6B161ACB1790CC66134A8CCA0D22A255ACB54A95055C9341B06694EB3D9AC952A14A24",
            INIT_RAM_05 => X"5CAE572B95C1D8EC76DA6D2E533B9ED2E9F6D60B8DC6F546B05D29D6CA9602EF26B0CC66",
            INIT_RAM_06 => X"0F37CB81C4F586C29EED37CB9988B25424950976D63B5FB3EA773D9EEFB7DBEDF6FB7DBE",
            INIT_RAM_07 => X"130B85CA653793D8A8172A241982E68A41201219BC9AC9138244680F1553C4EC501B14D8",
            INIT_RAM_08 => X"584A3C866114A93BAAF269553E47007BC85C5009BC920ACD844DAAD63A1D1622A850281C",
            INIT_RAM_09 => X"DF6FB7DBEDF6FB7DBE7D2E572B95CAE0EC761AED2E773DA6D36BA537AC05D2AD61BED46F",
            INIT_RAM_0A => X"0A2822111C56291C142F078B85E6FC813DDCB0C80B9984A8492B16CC170E1B5FB3EA7B3D",
            INIT_RAM_0B => X"952A358A8D1360ABDC910995026D66B75A2ED6CABC9E3944A5CEA6F22A2C266D166AB359",
            INIT_RAM_0C => X"586B35BECD60B8CC2F172A3B82D126A93D2A544A74561122564026F22A13DA291092C426",
            INIT_RAM_0D => X"2E48163F6FB3EE777CDF6FB7DBEDF6FB7DBE5CAE5F4B95CAE170761AED369B4DA4CA42B0",
            INIT_RAM_0E => X"0F4813D228CF723118F20702B5127053181591171BEDF704824120D1585BE1A8B6622C1A",
            INIT_RAM_0F => X"542A550A89509AC52A542A6552A54AA153DC5017B49225089952A8136B150A8700984CDF",
            INIT_RAM_10 => X"1A8D769B49927D602ED60B85DAC37EB151329519BC8A894D87C9295447B40A6D1257C8A8",
            INIT_RAM_11 => X"D14813C5C0D068B85C2E09163B53C3EE7B3DDF6FB7DBEDF6FB7DBE7D3E9F4FA5CAE17076",
            INIT_RAM_12 => X"EE5844DA4545843C240E66A51590F6AA3159CD5642A140A0309D9A8CE6BB8E07048B45A2",
            INIT_RAM_13 => X"952C05BACD16A85C2FD66B2D5ACF64A95266954AB596C136B04DAA951995226F2285C159",
            INIT_RAM_14 => X"7D3E9F4FA7D2E170761AED369B4742C0DE6F580BAE42E170BA5466D619BC866D519A53AC",
            INIT_RAM_15 => X"4C35FB961F248A41209137D3C5C2E068B81CCC66963B55CCEEF93D9EEFB7DBEDF6FB7DBE",
            INIT_RAM_16 => X"9169245A491691412291772C41EB1584BD9ACD566B3286C35DB0D8ACC81AFDBCA27AA552",
            INIT_RAM_17 => X"D66B26733DA0E3EE78FBCCD60B0371B85DECF61BC5BAC956B359ACD66B3596C54098D122",
            INIT_RAM_18 => X"DF6FB7DBEDF6FB7DBE9DBEA76FA5CAE4EC761ADCEE532372C163AC584C8DE2E957B05DAC",
            INIT_RAM_19 => X"6B955AEDF6BD493D0F88E4BB61E91381C1A29158A3C5C2E171BE1CC8A9A65B67D4EE7BBE",
            INIT_RAM_1A => X"745B2536C742A349A4912853CA05038349A45087A45629148940A04F07BB81C4F155AE96",
            INIT_RAM_1B => X"78AC05C6F37AC2653299BC5E333BA7DFEEB93C6DAE8F1782C0DC2E176B7596A54BA150A8",
            INIT_RAM_1C => X"276B267F67DCEE7B7CDF6FB7DBEDF6FB7DBE9DCEE76FA7D2E46C35B95C9E0F0372C160B0",
            INIT_RAM_1D => X"D2C8A456250075C0550A15428144F15427DCA954A33DC90380B8DF9048A3C5CCC173B516",
            INIT_RAM_1E => X"DA4CE673258CC962B0780BB5BAC955B254A854CA84DE4D2F9349E4D26974BA412E904C26",
            INIT_RAM_1F => X"B93C1E06E170B8DEB0381C0E0B0381C162B0582C16070382C265B41BAE4F1B6DB6D369B4",
            INIT_RAM_20 => X"6FA7AB398CC660248D0A6B267F77D4EE7B3DDF6FB7DBEDF6FB7DBE9DCEE76FA7D2E46B73",
            INIT_RAM_21 => X"54CAA54A9541A04CA99509B4826F2489419A8C053A8A688156A59288139AF1991489BEDF",
            INIT_RAM_22 => X"788DCF0B97DCED72B95C9E0F0383C0DBEFB6BA3C56270179BC5FAD17EB7592AD66B2532A",
            INIT_RAM_23 => X"9DCEEF8FA7D2E46DB4B93C1E02D169B8DC70381C16070382C0E070589C0E070381C0DC6F",
            INIT_RAM_24 => X"0A64A44985028140DF0E27835168B04A2C95CC7B266377D5F27B3DDF6FB7DBEDF6FB7DBE",
            INIT_RAM_25 => X"582C5622F178BC5E2F178BF59ACB64A9D0A9952A0CDE47409B48A690072B2149064AB352",
            INIT_RAM_26 => X"B94C9E2F0783C5E0F058CCB6CB97DBEA76FA9DBEDF4B95C9E07037FBCCE673358CC962B1",
            INIT_RAM_27 => X"DF6FB7DBEDF6FB7DBEBE4EE773B9DBE8EC76B95CAE572783C26532994CA653299CCE66F1",
            INIT_RAM_28 => X"D2488BD9A4B5662194880521F925048AC49E2E37CB9988B45A2D98CD6B5E4377DCF67B7C",
            INIT_RAM_29 => X"3C0E3EFF7DAED66B339ACCE673399CCA66B1589C0DE2E16EB75B2AD62A652A9741984C66",
            INIT_RAM_2A => X"FB6D7EDB5FB6D3EDB4FB6DB69B5DA6D369B4DA5CEE9B51BAE5F73B9DCEDF6B95CAE57278",
            INIT_RAM_2B => X"0E6B1E4787DDF27B3DDF6FB7DBEDF6FB7DBEBE5F2777C9DBE970761A8D46BB4DA5CF6DB6",
            INIT_RAM_2C => X"D6EB2552A954AA54A833792C4DFEE461BF108864A21105048A449ED1489BE5C8B35E319A",
            INIT_RAM_2D => X"7DBEE76FA7DBEDF4FA7D2E572381C7DFEFF7FBFDF6DB6BA5D2673399CCD62B1589BC5E6F",
            INIT_RAM_2E => X"3B1D8EC363B0D8F0373C0DC6E781C0E070781B1E06C781B0E06E361BFDBEDF6FB0DCF0B9",
            INIT_RAM_2F => X"B1589401CEA660385C903A266377DDF27BBEDF6FB7DBEDF6FB7DBEBE5F2F97C9DCED7276",
            INIT_RAM_30 => X"DACD6673358AC4E1AD170BC5DADD60BA552A545A84DA26FF712DDCA9238299250B81C0A0",
            INIT_RAM_31 => X"5CAE4F0373C1E0F0781C1E172B97D2E5F4FA7D2E572FA5C9E0F0783C1E06E37FBEDBEFB6",
            INIT_RAM_32 => X"BE5F2F93B9DBE972B83B1D8EC763C1E0F0783C1E0F0785C9E172B95C2E572B95CAE172B9",
            INIT_RAM_33 => X"2AD491D920EC8244E0B169140D74AB7CB8DF0E4A5E6377DDF27B7CDF6FB7DBEDF6FB7DBE",
            INIT_RAM_34 => X"7D3E972781C1E0F0381C7DF6DB59ACCE6A2F78BC160B0170B759AC543A35824B0B7C3918",
            INIT_RAM_35 => X"5CAE572B95CAE572B97D2E572783C1E0F0785C9E0F0781C0E0F0785CAE572B97D3E9F6FA",
            INIT_RAM_36 => X"DF6FB7DBEDF6FB7DBEBE5F2F97CBE5F1F4B85C1D8F0783C1E172783C2E4F0785CAE572B9",
            INIT_RAM_37 => X"D64A9D12812585BFDC4B750290F8C87B4BA4D1689C0D86C76BB49E6F89A66787D5F37D3D",
            INIT_RAM_38 => X"3C0E0F0785CBE972FB5CBEDF4FA5CAE572B93C0E071F7DB6DB6933DA5CE6732581BD61AC",
            INIT_RAM_39 => X"5C9E0F0B95CAE172B97D2E572FA5CAE5F4B95CAE572B93C1E0F0B95CAE5F4B93C1E0F038",
            INIT_RAM_3A => X"90791E2787DCF77D3DDF6FB7DBEDF6FB7DBEBE5F2F97CBE3E972B85C2E0EC783C1E0F078",
            INIT_RAM_3B => X"FBEDB6BB49AAC562F0176B1506694692405CACA5B25524B58B4826D2690381C0E37DBEDF",
            INIT_RAM_3C => X"5CAE572FA5CAE572B95C8E070381C1E070B95CAE572FB7D3ED72FB5CAE572781C0E06FF7",
            INIT_RAM_3D => X"5C1D970783C1E0F0783C1E172787D2E572B95CAE572B95CBE972B97D2E572FA3C1E17278",
            INIT_RAM_3E => X"D2792C5A22E27838DF2E791E2387DCF6F9BEDF6FB7DBEDF6FB7DBEBE5F2F97CBE4EDF4B8",
            INIT_RAM_3F => X"7DBE972FA5CAE4F0783C0E3EFF7FBCD666B1580B7592A532A344DF0E360AA96EE48B4BA4"
        )
        port map (
            DO => promx9_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_13,
            RESET => reset,
            AD => promx9_inst_6_AD_i
        );

    promx9_inst_7: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"5CAE572B93C1E172785CAE5F4FA7D2E572B95CAE4F0781C0E071F7FB8E070785CAE572FA",
            INIT_RAM_01 => X"BE5F2F97CBE4EDF4B85C1D8F0783C1E172785C9E0F0B95C1E172B95C3E972B85CAE570B9",
            INIT_RAM_02 => X"4F5652C14ACA8349A4F2793C9A4F2382C361D109A66389DCF6F93DDF6FB7DBEDF6FB7DBE",
            INIT_RAM_03 => X"FBFDF6DB5DB6DB6DB4FB8E0F0383C2E572B91C3E8F0783C0DF6DB5999C05D6A741984920",
            INIT_RAM_04 => X"5C1E170785C1E0F0783C2E570B93C1E0F0B97D2E572FA5CAE4F0783C2E572B93C1E0F037",
            INIT_RAM_05 => X"DF6FB7DBEDF6FB7DBEBE5F2F97CBE5F1F4B83B1D8EC381C1E0F0783C2E0F0783C1E0F078",
            INIT_RAM_06 => X"DB6D2646FF64A94D61F1F723118EE0784DA4916904C261319848E0112A562377DCF77DBE",
            INIT_RAM_07 => X"1B8DD72785CAE4F0381C7DFEDB6DB6DB6D74DA4D6E97499CCEE8381C2E4F0B95C8E071F7",
            INIT_RAM_08 => X"1B8E0F0383C1E070783C0E0F0363C1D8F0783C1E0F0B83C2E4F0B95CAE5F4B95C9E0F037",
            INIT_RAM_09 => X"131A266789DDF27BBEDF6FB7DBEDF6FB7DBEBE5F2F97CBE5F170B85C1D86C371B8E06E36",
            INIT_RAM_0A => X"373C265B51B8DC6E381BFDF6933587B2D464B0C8335180E693C826D1098CC24D1071C024",
            INIT_RAM_0B => X"5CAE5F4FA5CAE4F037FB0DC6E781C2E572383C0E3EDB61B6DB6DB6DA5D369B4BA5CA66F1",
            INIT_RAM_0C => X"3B1D8EC371B0E06E381B8E0F0381C1E0F0783C1E0EC781C0E0F0783C2E4F0B93C1E0F0B9",
            INIT_RAM_0D => X"3369749610EE4AA41ECE67266377DCF67BBEDF6FB7DBEDF6FB7DBEBE5F2F97CBE5F1F4B8",
            INIT_RAM_0E => X"DA6D66772BA5CAE933784C9E0B0378B96133DAEDB6D3599BC45D2A12488385C915884C66",
            INIT_RAM_0F => X"5C9E0F0783C1E172B95CAE572B95C9E0F0781B8DC6E371B9E172385C9E071F7DB7DF6DB6",
            INIT_RAM_10 => X"BE5F2F97CBE4EDF4B85C1D970783C0E0F0783C1E0F0783C1E0F0783C1E0F0783C1E17078",
            INIT_RAM_11 => X"95092405ED20995226F238244A00F4409C4EA946562789DDF27BBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_12 => X"3C1E0F0781C7DFEFF7DA6DAE97499DD2E77378CCA6532782C05DACD56B0DD3399CCD622E",
            INIT_RAM_13 => X"5CBE972B95CAE572B93C2E572B93C1E0F0785CAE572B95CAE4F0783C1E070781B9E0F078",
            INIT_RAM_14 => X"DF6FB7DBEDF6FB7DBEBE5F2F97CBE5F1F4B85C2E0EC783C1E0F0B93C2E572B95CAE572B9",
            INIT_RAM_15 => X"376AA5128172C562B0385A8492090999522613696C5A4EE56735185069162789DCF77DBE",
            INIT_RAM_16 => X"3C0DC6E781B9E06E371C0DCF0373C1E0F1F6FBEDAE9B6BA4CE6733994CE6732994C9606F",
            INIT_RAM_17 => X"5C9E0F0783C1E1F4B95CAE4F0B95CAE572B95CAE4F0B93C2E572785C9E172B95C9E0F078",
            INIT_RAM_18 => X"D209562789DCF67BBEDF6FB7DBEDF6FB7DBEBE5F2F97CBE4ED70B85C2E170783C2E57278",
            INIT_RAM_19 => X"994CA653258AC160B0378BB592873EA85C7037EB5D026130995226132A44C261348A4562",
            INIT_RAM_1A => X"1C0E06C371B8DC6E37FB0DC6FF6FB7DBEFF6FB7DBEDB6FB7D86E781C7DF6DB5DB5D2E933",
            INIT_RAM_1B => X"5C1D8EC383C0E0F0783C1E0F0783C1E070783C1E0F0783C1E0F0783C1E0F0781B8DC7038",
            INIT_RAM_1C => X"334AA552A53092C41ED2CA85E789DCF77DBEDF6FB7DBEDF6FB7DBEBE5F2F97CBE5F1F4B8",
            INIT_RAM_1D => X"1B8E06E37FBEDAE93399CCA64B0582C160B0582C0DDEC9489251EC170BF58A9130984C26",
            INIT_RAM_1E => X"1A8D46A351AFD86BB41AED86BB61AED369B4DA6D369B4DA6D369B4DA6D26733BA5D2E9F6",
            INIT_RAM_1F => X"BE5F2F93B9DBE970B85C1D86DF71B7DFEE37FBFDC6FF7FB7DBEC361B0D86C361B0D86C36",
            INIT_RAM_20 => X"B57B3596A546974826954AAD4A954A9BC722F24935A789EDF27BBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_21 => X"783C5E0F0783C160B199ED070381C0DFEFB5DA4CE66B0582C560B0582C1606E174A048E6",
            INIT_RAM_22 => X"DA6D369B4DA6D36973DA5CEE773B95CEE772B95CEE572B94CEE532993C66532783C5E2F0",
            INIT_RAM_23 => X"DF6FB7DBEDF6FB7DBE7D3E9F53B7D5F170B81B0DB69B4DA5CF6973DA6D369B4B9ED369B4",
            INIT_RAM_24 => X"582C0DC6E378BBD422946B3D9ACB609A45A454CAA55625097B49E34F8775AB99ECF77DBE",
            INIT_RAM_25 => X"58AC160B0582C560B0582C1606F381BCDE7037BC3EEB93C0E06FF7DB6DA6732582C160B0",
            INIT_RAM_26 => X"995CA6532995CAE572B9DCEE772B9DCAE572994CA6532994CA64F0994CA64B078AC160B0",
            INIT_RAM_27 => X"344A45EB99DCF77DBEDF6FB7DBEDF6FB7DBE5CBE9F4FA7D2E570761B6D2E97399CCA6532",
            INIT_RAM_28 => X"FBEDA6B73992C162B0582C0DC6E371BBD8E7125AB59ECD62A349A4D2CA654E81379049A4",
            INIT_RAM_29 => X"994CA64B058AC160B0582C160B0582C160B0382C1606E379C1606E371BB6A785CAE57278",
            INIT_RAM_2A => X"1B6D2E733B94CA6532995CA6532994CA6532B95CEE772B94CAE532B94CA6532994C9E132",
            INIT_RAM_2B => X"D25884D2A954AA556AD60BD62B9BE4F67BBEDF6FB7DBEDF6FB7DBE5CAE572B95CAE57078",
            INIT_RAM_2C => X"582C2E8373C2E572781C0E3EFB6DA5CA66B1582C1606F371B85DAC944A355AC16EB153A5",
            INIT_RAM_2D => X"B9DCEE773B9DCEE733B94CEE533995CA6532994CA6532994CA64F178BC5E0F058AC1E0B0",
            INIT_RAM_2E => X"3C0E0F0B85CAE17238FB6DB6974DA5CB6974DA5D2E973BA6D369B4DA6D369B4DA6D2E774",
            INIT_RAM_2F => X"F629AD5ACD66B6542691489412250E91512AD60BD62FA9ECF77DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_30 => X"DA6D36973DA5CEE572BA4CEE9B6FBAE572B95C9E0F038FBEDB6932582C160B0581B8DC6E",
            INIT_RAM_31 => X"1B0D46A361A8D46A351AED06BB41AED06A35DA6DB6DB4DA6DB69B4DA6D369B4DA6D369B4",
            INIT_RAM_32 => X"DF6FB7DBEDF6FB7DBE3C2E4F0B95CAE4F0B83C0D86DF6FB8D76C351AFD86BF61B0DBEC35",
            INIT_RAM_33 => X"9ABC5E0B0582C0DE6F37EB2D5ACD68B75929D2488BCE00E07AB3A4B60BE66FA9EDF37DBE",
            INIT_RAM_34 => X"1B8DC6DF6FBFD86C361B7D86A35DB6D86BB6DB6DBEDF6FB8E0F0785CAE572B91C1E3EFB5",
            INIT_RAM_35 => X"3C1E0F0781C1E0F0783C1E0F0783B0E070381B0D8EC363B0DCEC371B0D8EC371C0DC6E36",
            INIT_RAM_36 => X"B62C66AFBBE4F77DBEDF6FB7DBEDF6FB7DBE5CAE5F4FA5CAE572B95C9E172783C1E0F078",
            INIT_RAM_37 => X"FB9E3EE785C9E0F038DB5D264B0582C1606F378BA55ACD66B45B6A13480BC1CEE0783BA4",
            INIT_RAM_38 => X"3C1E0F0783C1E0F0783C1E0F0783C0E070371B8DC70361B8DC6E371BFD86FF6FBFDC6E38",
            INIT_RAM_39 => X"5CAE572B95C1E172B93C2E572B95C9E172B95CAE572B95CAE570B93C2E4F0B83C1E0F078",
            INIT_RAM_3A => X"54C88BDDCEE77141A5D62C66AFA9ECF77DBEDF6FB7DBEDF6FB7DBE7D3E972FA5CBE972B9",
            INIT_RAM_3B => X"1B8DC6FB6DB6DB6BB6FB8E3EFB5FB9E172B93C7DEE932992C5606F378BB59AC168B45DEC",
            INIT_RAM_3C => X"5CAE0F0783C2E572785C9E0F0783C1E0F0783C1E06E783C0DCF0783C1E06E371B8DC6E37",
            INIT_RAM_3D => X"5CAE5F4FA5CBE972B95CBE8F0B95CAE572B83C3E972B95CAE572B95CAE572B95CAE572B9",
            INIT_RAM_3E => X"582C05D6AD60B8E02F95691BE1C0E286446817CCFED3B9EDF37DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_3F => X"3C1E06E371B8DC6E371B8DC6FB599AC667F71C0E36B35FB8E0F0B93C1E071B499CC9E2F0"
        )
        port map (
            DO => promx9_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_15,
            RESET => reset,
            AD => promx9_inst_7_AD_i
        );

    promx9_inst_8: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"E7F1F8DC6E36DB4D9EC2DB6CB549A40DC6A26940EABB6DB71F9FD7F3FBFCFF7FBFDFEFF7",
            INIT_RAM_01 => X"EFF5FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FBFE7F3F5FBFDFEFF5F9FD7",
            INIT_RAM_02 => X"EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEBF7FAFDFEBF7FAFD7EBF5FAFD7EBF7FCFDF",
            INIT_RAM_03 => X"F3F9FEFF7FBFDFEFF7E7F3F9FDFE7F7F9FCFE7EFB7DBEDB6FB7DC6E373F9FDFEFF7FBFDF",
            INIT_RAM_04 => X"F3F5FBFD7EFF3F9FCFE7F1B8DB6DB69B1D8DB6D96A93C81B8D44916140E9BA6DB71F9FD7",
            INIT_RAM_05 => X"EBF5F9FD7EBF9FCFE7F3F9FDFE7F3F9FDFE7F3F9FCFE7F7F9FCFE7F7F9FCFE7F3F9FCFE7",
            INIT_RAM_06 => X"E373F9FCFEFF7FBFDFEFF7FBFDFEFF7FAFDFEFF5FAFD7EFF5FBFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_07 => X"5938E9B96DB71F9FD7F3F9FCFF7FBFDFEFF7E7F5FAFDFEFF7F9FCFE36FB7DAED76FB7DBE",
            INIT_RAM_08 => X"F3F9FCFE7F3F9FCFE7EFF5FAFD7E7F3F9DC7E771B6DB6CB65AEB65A6D36690B69244A071",
            INIT_RAM_09 => X"EBF5FAFD7EBF5FAFCFE7F3FBFE7F3F9FCFE7F7F9FDFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7",
            INIT_RAM_0A => X"E36FB7DAED76BB6DBEDF71B9FCFE7F7FBFDFEFF7FBFDFEFF7F9FD7EFF3F9FCFE7F5FAFD7",
            INIT_RAM_0B => X"A2491F6B23892080714938E898EDB71B9FD7F3F9FEFF7FBFDFEFF7EFF5FAFDFEFF7FBFCF",
            INIT_RAM_0C => X"F3FBFCFE7F3F9FCFE7F3F9FCFDFF3F7FAFD7EBF3F9FCFE7F1B8DC6E36DB6DA6C2DD6CB54",
            INIT_RAM_0D => X"E7F3F8FCFE7F3F9FCFEFF5FAFD7EBF3F8FC7EBF5FAFE7F3F9FDFE7F7F9FDFE7F3F9FCFEF",
            INIT_RAM_0E => X"EFF5FBFDFEBF7FAFCFE36FB5DAED76BB5DBEDF71B8DCFE7F3FBFCFEFF7FBFCFE7F3F9FCF",
            INIT_RAM_0F => X"DB69B2D6DAAD12691371B28E23818080606144B8E8985DB71B9FDFF3FBFEFF7FBFDFEFF7",
            INIT_RAM_10 => X"F7FBFCFEFF3F9FCFE7F3F9FCFE7F3F9FCFDFEFF9FBFE7EFF7FAFD7E7F7F9DCEE771B8DB6",
            INIT_RAM_11 => X"E7F3F9FDFE7F3F9FCFE7F3F9FCFE373F8FCFE7F3F9FCFEBF1F8FD7EBF9FDFE7F7F9FDFEF",
            INIT_RAM_12 => X"F3FBFEFF7FBFDFEFF7EFF7FBFDFEFF7FBFDFE36FB7DAED76BB5DBEDF71B8DCFE7F3F9FCF",
            INIT_RAM_13 => X"E773B9DB6DB6DB4DA6CF59606F3692C93481240C040180C080405044B4E8975DB6DB9FD7",
            INIT_RAM_14 => X"F3F9FCFE7F7FBFDFEFF3F9FCFE7F3F9FCFE7F3F9FCFE7EFF7FAFD7EBF7FBFDFEBF7FBFCF",
            INIT_RAM_15 => X"DB6FB8DCFE7F3F9FCFE7F3F9FC6E7F3F9FCFE371B8DC6E371B7DC6E371B8DC6E373F9FE7",
            INIT_RAM_16 => X"38B8E6985DB71B8FD7F3F9FEFF7FBFDFEFF7EFF7FBFDFEFF7FBFCFE7F1B7DAED769B4DBE",
            INIT_RAM_17 => X"E7F3F9FCEE3F3B9DC6DB6DB2D9EC2D9689135098460302014060201006030180C0604048",
            INIT_RAM_18 => X"D76BB4DAEE377FCFE7F3FBFCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FBFDFEFF7FBFDF",
            INIT_RAM_19 => X"E7EFB5DAECF67B4DA6D76BB7DB6DF6FB7DBEDF6FB7DBEDF6DB7DAEDF6BB5DAED369B4DAE",
            INIT_RAM_1A => X"1406030180C060303830B8E598EDB6DB9FD7F3FBFCFF7FBFDFEFF7F3F7FBFE7EFF7FBFDF",
            INIT_RAM_1B => X"EFF7FBFCFEFF3F9DCEE371B8DB6DB69B4D9EAAB8D1240241004020101206018181008020",
            INIT_RAM_1C => X"CB65B2D95C76170B85C2E172DB6EFF9FCFEFF3FBFCFE7F3F9FCFE7F3F9FCFE7F3F5FBFDF",
            INIT_RAM_1D => X"EFF7FCFE7EFF7FBFDFE36FB4DA6D36572D9ECF65B4DA6D369B5DA6D369B4D96CB67B3D9E",
            INIT_RAM_1E => X"1008070181408060201008030180C060303028B8E5985DB71B8FD7F3F9FEFF7FBFDFEFF7",
            INIT_RAM_1F => X"EFF7FBFDFEFF5F9FCFE7F3B9DC6DB6DB5DA6CF6166892449406030180804018181004020",
            INIT_RAM_20 => X"C763B1D8EC2E170B85C2DD6EB6DB6D96CB65B2E3B8DE7F3F9FCFE7F3F9FBFE7F3F9FBFE7",
            INIT_RAM_21 => X"F3F9FCFF7FBFDFEFF7F3F9FCFE7F3F7FBFDFDF6FB4D9DC6E170B85C6E3B1D96CB65B2D8E",
            INIT_RAM_22 => X"180804018100C040201008060201808040300C08030180C060302828B8E598EDB6DB9FD7",
            INIT_RAM_23 => X"EFF7FBFD7EFF7FBFDFEFF3FBFCFE371B6DC6D367B2B5469AA8A050308C06018100806030",
            INIT_RAM_24 => X"C763B1D96CB65B2D96C765B1D85C2E170B75BAE16EB6DB6DB6CB6DC771BCFE7F3F9FCFE7",
            INIT_RAM_25 => X"28B8E6996DB6DB8FD7F3FBFCFF7FBFDFEFF7F3F9FCFE7F3F9FBFDFDF6FB4DA6D36170B8D",
            INIT_RAM_26 => X"280E040200C0604030200C06018100E050201006060201C0806038100604020100804028",
            INIT_RAM_27 => X"E3F7FAFE7EFF7FBFDFEFF7FAFCFEFF3F9DCFE771B7DB6D76BB4D9ECADD6AAAA140C04038",
            INIT_RAM_28 => X"EFEFB5D9ED367B3D9ECF69B4DA6D369B4DA6D369B4DA6CB65B1D8EC763B0B95C2E16EB96",
            INIT_RAM_29 => X"0C060302008080203828BCE6996DB6DB8FD7F3F9FDFF7FBFDFEFF7F7F9FDFE7F3F9FBFDF",
            INIT_RAM_2A => X"C6DD6A8D21008060302010060201006040381810080301810060201408070201C0806040",
            INIT_RAM_2B => X"D769B4DA6CB69B4DD7EBF1FAFDFEFF3B8DC6E371B6DB6DF6FB6DC6E36DB7DB6D769B3D96",
            INIT_RAM_2C => X"F3F9FCFE7F3F9FBFDFE7F3F7DBED76BB6DB6DF6FB7DBEDF6FB7DBEDB6FB7DB6DB6BB6DAE",
            INIT_RAM_2D => X"20080702018080604010060302014060402028C0E9BA6D36DB8FD7EFF9FCFF7FBFDFEFF7",
            INIT_RAM_2E => X"DF6DB6DB6D769B3D85C2DB6A903200C04030200E050280C0806020180C080401C100A040",
            INIT_RAM_2F => X"E7F3FAFCFE7F3F9FCFE373F9FBEDF71BAFDFE7F1B7DBEDF6FB7DB6DF6DB7DBEDF6FB7DBE",
            INIT_RAM_30 => X"EBF9FEFF7FBFDFEFF7F7F9FCFE7F3F9FCFDFEFF7FBFCFE371B8DCEE7F3F9FDFE7F7F9FD7",
            INIT_RAM_31 => X"1C1008040200E08040200C08030180C060301008040200C060302830C0F0BA6DB71B9FD7",
            INIT_RAM_32 => X"DF6DB7DB6DB6DB6DB6DB6DB5DAED769B2D8DC2D968903308806040201006020100606040",
            INIT_RAM_33 => X"EBF7FAFD7EFF5FBFD7EFF5FBFD7EFF5FAFDFEFF3F9FCFE3F5FAFC7E371B7DBEDB6FB6DBE",
            INIT_RAM_34 => X"494B32DB6DB6DB8FD7EFF9FCFF7FBFDFEFF7F3F9FCFEFF3F9FCFE7EFF7FBFCFE7F3F9FCF",
            INIT_RAM_35 => X"181007038180804028201009040200E0805018100A0301C0C06030100A040100C0803028",
            INIT_RAM_36 => X"E771B7DBEDF6FB6DBEDB6FB6DBEDB6DB6DBEDB6DB5DAED367B2D85BAD968913448804040",
            INIT_RAM_37 => X"EFF7FBFDFEBF3F9FD7E7F5FBFD7EFF7FBFDFEFF7FBFDFEFF7FAFD7EFF5FAFD7E7F5FAFDF",
            INIT_RAM_38 => X"140C04018100A04028695D72DB6D371B9FD7EFF9FEFF7FBFDFEFF7F7F9FDFE7F7F9FCFE7",
            INIT_RAM_39 => X"BAD966913550808048180C060401C10080201C1007040201008048241008040201006030",
            INIT_RAM_3A => X"EBF7FAFD7E7F7FCFD7E7F1B7DB6DB6DB6DAEDB6DB6DB6DB6DB6DAED76BB5DA6CF67B2B7D",
            INIT_RAM_3B => X"F3F9FCFE7F7F9FDFE7EFF7F9FD7E3F3FAFD7E7F7FAFDFEFF7FBFDFEBF7FBFD7EFF5FBFDF",
            INIT_RAM_3C => X"2810070402410070301C0E040200C080303081E5B4DA6DB71B9FCFEBF9FCFF7FBFDFEFF7",
            INIT_RAM_3D => X"D769B5DA6CF65B0B85B6D568913490805040200C06030241446040201008030201008050",
            INIT_RAM_3E => X"EBF7FBFDFEFF7FBFDFEFF7FBFD7EBF5FCFD7E7F5F9FC7E371B7DBEDB6DB6DB6DF6DB5DAE",
            INIT_RAM_3F => X"EBF9FCFF7FBFDFEFF7F7FBFDFE7F7F9FCFE7EFF7FBFD7EBF1FAFD7EBF5FAFD7EFF5FBFDF"
        )
        port map (
            DO => promx9_inst_8_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => promx9_inst_8_AD_i
        );

    promx9_inst_9: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"18100804018184A048281009030200E08030201204010100A050599665B4DB6DB6DB9FD7",
            INIT_RAM_01 => X"E36DB6DB6DB6BB6DAED369B4D9ECB6570B75B6D5669135508040301C1206030201408030",
            INIT_RAM_02 => X"EBF5F9FD7EFF7FBFDFEBF7FBFD7EFF5FBFDFEFF7FBFD7EBF9FCFD7EFF7FBFCFEBF3F8DC6",
            INIT_RAM_03 => X"BAE5B4DA6DB6DB9FD7EFF9FCFF7FBFDFEFF7F3F9FCFE7F7F9FDFE7EFF7FAFCFEBF3FAFCF",
            INIT_RAM_04 => X"1C0E080302014480381C10090381C184C24828100C2401C0C08038181404018140805061",
            INIT_RAM_05 => X"EBF5FAFCFEBF3F9FCFE771B8DBEDB6DB6DAED769B4D9ECB616EB75B2D326913448804030",
            INIT_RAM_06 => X"EFF7FAFCFEBF3FAFD7E7F5FAFD7EBF5FBFDFEBF7FBFDFEFF7FAFDFEFF7FAFCFEBF9FCFD7",
            INIT_RAM_07 => X"1C10040181008050F3C767B3DA6DB6DB9FD7EFF9FCFF7FBFDFEFF7F7FBFDFEFF7F9FCFE7",
            INIT_RAM_08 => X"B2D125913388804040140C0803820140A24820120A03820144A24020100A0501C0807040",
            INIT_RAM_09 => X"EFF7FAFD7EFF9FCFD7EBF7FAFD7EBF5FBFD7EBF3F8DC7E371B6DB6D769B3D9ECB616FB65",
            INIT_RAM_0A => X"F7FBFDFEFF3F9FCFE7EFF7FBFD7EBF3FAFC7EBF5FAFD7EBF5FBFDFEFF7FBFD7EFF5FBFDF",
            INIT_RAM_0B => X"200E080511C0C080401C0E0402814060614CC2E9B4D9EDB71B9FD7F3F9FCFF7FBFDFEFF7",
            INIT_RAM_0C => X"DF6DB4D96C6E16EB75AAD126903240E0402828080804020144A25028920A04028920A050",
            INIT_RAM_0D => X"EBF7FBFDFEFF7FBFDFEFF7FBFD7EBF9FCFD7EFF5FAFD7EBF5FBFD7EFF5FAFCFE3F1F9DB6",
            INIT_RAM_0E => X"EFF9FCFF7FBFDFEFF7F3FBFCFEFF3FBFCFE7EFF5FBFD7EBF5FAFD7EBF5FAFD7EBF5FBFDF",
            INIT_RAM_0F => X"281408061281008050240E08050180E0804018120702018060B38ECB67B3DA6D371B8FD7",
            INIT_RAM_10 => X"EBF7FAFD7E7F3F9FC6DB6DB4DA6C7616EB65AA51258F3200A06020140A07048201008050",
            INIT_RAM_11 => X"EBF5FAFD7EBF5FAFDFEFF7FBFD7EFF7FBFDFEFF7FAFD7EBF9FBFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_12 => X"CB65B2DA6DB6DB9FD7EFFBFCFF7FBFDFEFF7F7FBFDFE7F3F9FCFE7EFF7FBFD7EBF5F9FC7",
            INIT_RAM_13 => X"100A04040240E08048201208050309009059281008051280E0A0401C0C0702818081558E",
            INIT_RAM_14 => X"EBF5F9FD7EBF7FAFD7EBF5FAFD7EBF3F9DC6E36DB4D9EC7616EB65AA4D268D3100804020",
            INIT_RAM_15 => X"EFF7FBFD7E7F5FAFD7EBF5FAFD7EBF5FAFDFEBF7FAFDFEFF5FBFDFEFF7FBFD7EFF9FAFDF",
            INIT_RAM_16 => X"200C060281C0E12585CB65B2DA6DB71B8FD7EFF9FEFF7FBFDFEFF7F7F9FCFEFF3FBFCFE7",
            INIT_RAM_17 => X"AA4D2289210080402010080503028120804024184A05128900A251288E07040240E08040",
            INIT_RAM_18 => X"EFF7FAFDFEBF5FBFDFEBF7FAFD7EFF5FAFD7EFF7FBFDFEBF1F8FC6E36DB5DA6CB616EB55",
            INIT_RAM_19 => X"F3F9FCFE7F3FBFCFE7EFF7FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFDFEBF7FBFDFEFF5FBFDF",
            INIT_RAM_1A => X"288E09048281007040240C05038180C16575CB67B3D96DB71F9FD7EFF9FDFF7FBFDFEFF7",
            INIT_RAM_1B => X"DF6DB5DA6C7616DB55A24D226611C100502018080504820100703018100805128900A250",
            INIT_RAM_1C => X"EBF7FBFDFEFF5FBFDFEFF7FBFDFEBF5FBFCFEBF7FBFCFE7F7F9FD7E7F7F9FCFE7F1F9FC6",
            INIT_RAM_1D => X"EFF9FCFF7FBFDFEFF7F3F9FDFE7F3F9FCFE7EFF7FBFD7EBF5FAFD7EBF5FAFD7EBF5FAFDF",
            INIT_RAM_1E => X"180C0805028900906128900A240241006028200804038140E1A775CB65B2D9EDB6DBAFD7",
            INIT_RAM_1F => X"EFF3F8FCEE371F9FC6DB6DB4D9ECAE16DB65A24B1E620100E07028180C05048241008030",
            INIT_RAM_20 => X"EBF5FAFD7EBF5FAFDFEFF7FBFDFEFF7FBFDFEFF7FBFD7EBF5FAFD7E7F3F9FCFE7F3F9FDF",
            INIT_RAM_21 => X"CB65B2DA6DB71F9FD7F3F9FCFF7FBFDFEFF7F3F9FDFE7F3F9FCFE7EBF7FAFD7EBF5FAFD7",
            INIT_RAM_22 => X"140E07040280E080401C0C0A24830920905028920A040280E040381C0C04030140E18575",
            INIT_RAM_23 => X"E7F1F9FCEE3F3B9DC6E371B8DCFE371B8DB6DB6DB4D96C6E16CB55A24B18420100805030",
            INIT_RAM_24 => X"EBF7FAFD7EBF5FAFD7EBF5FAFD7EBF7FBFD7EFF7FBFDFEBF7FAFDFEFF7FBFDFEFF5FAFDF",
            INIT_RAM_25 => X"1C0804028180816575CB65B2D9EDB6DB9FD7EFF9FDFF7FBFDFEFF7F3F9FCFE7F3F9FCFDF",
            INIT_RAM_26 => X"9A49112301C0C03020100A04030241008038200C08040309409051241208040280E07048",
            INIT_RAM_27 => X"EFF7FBFD7EBF5FAFDFE771F9FC6E371F9FC6DB71B8DB6E371B8DB6DB6DB4D9EC2DD6CB55",
            INIT_RAM_28 => X"F3F9FBFE7F3F9FCFD7EBF7FAFD7EBF5FAFD7EBF5FAFD7EBF5FBFDFEFF7FBFD7EFF7FBFDF",
            INIT_RAM_29 => X"28900803020100705114080402018080C36DCB65B2D96DB71F9FD7EFF9FCFF7FBFDFEFF7",
            INIT_RAM_2A => X"DB69B4D9EC2DD6DB55A240CC240200C08020100807048181009038281009050281208051",
            INIT_RAM_2B => X"EBF7FBFDFEBF7FAFDFEFF7FBFDFEFF7F9FCFE3F3F8DC6E371B7DBEDF6DB6DB6DF71B8DB6",
            INIT_RAM_2C => X"F3F9FDFF7FBFDFEFF7EBF5FAFD7F3F5FBFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_2D => X"289209050200E060503090060301C0E0704018080702014080A36DCB65B2D9EDB6DB9FD7",
            INIT_RAM_2E => X"DB6DB5DB6E371B6DBEDB69B4D9EC75D6EB549A38C90401C1008028100807040280E08040",
            INIT_RAM_2F => X"EBF5FAFD7EBF5FAFD7EFF5FBFD7EFF7FBFDFEFF7FBFDFEBF5F9FCFE771B6DB6DF6DB6DB6",
            INIT_RAM_30 => X"BAE5B2D9EDB6DB9FD7F3FBFCFF7FBFDFEFF7EBF5FBFD7EFF5FBFD7EFF5FAFD7EBF5FAFD7",
            INIT_RAM_31 => X"1C140502028900903020144C250200C060503090070401C0C06030140804020100A0916D",
            INIT_RAM_32 => X"E371B8DB6DB6DB7DAED76DB6DBEE371B8DB6DB69B4D9ECB616DB559A2486040180806030",
            INIT_RAM_33 => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFDFEBF5FBFD7EFF7FAFDFEFF7FBFDFEFF3F9FCE",
            INIT_RAM_34 => X"240C05038100C0711CBAE5B2D9EDB71B9FD7EFF9FDFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_35 => X"921C44020180C060401C0E0902018140903024100E250240E0A0512C8E05030140E06038",
            INIT_RAM_36 => X"EFF5FBFE7EBF3FAFCEE371B7DB6D76DB6DAED36DB6DC6E771B8DC6DB6DB4D9ECB616CB55",
            INIT_RAM_37 => X"EBF7FAFDFEBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFDFEFF7FBFDFEFF7FAFDF",
            INIT_RAM_38 => X"1C0E0604820144C26128984A2302016480D3B6E5B2D96DB71B8FD7F3F9FCFF7FBFDFEFF7",
            INIT_RAM_39 => X"DB69B4D96C2DD6AB347990050200C0C060401C0808040140E0806120144E250281008048",
            INIT_RAM_3A => X"EBF5FBFD7EFF7FBFDFEFF5FCFD7EBF5F8FC6E371B6DBEDB6BB5DAED76DB8DC7E371B6DB6",
            INIT_RAM_3B => X"F3F9FDFF7FBFDFEFF7EBF5FBFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_3C => X"24120C250288E0A03020120904044A25248949224C251181848092A6E172D96D371B8FD7",
            INIT_RAM_3D => X"DB71B8DCFE36DB7DB6D769B3D96C2DD6A934490A07038180C06028289007051200C0A248",
            INIT_RAM_3E => X"EBF5FAFD7E7F3F9FCFEBF5FAFD7EBF7FAFDFEBF7FAFDFEFF3F8DCEE371B7DB6D76BB4DA6",
            INIT_RAM_3F => X"8A5D72D96D36DB9FD7F3F9FCFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7"
        )
        port map (
            DO => promx9_inst_9_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => promx9_inst_9_AD_i
        );

    promx9_inst_10: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"14144905128920905124120A048240C0603030A2512924934954AA69AC9247128944A271",
            INIT_RAM_01 => X"E771B7DB6DB6BB6DB6E371B8DC6E371B6DB6D367B0B85BAD568913200A050381C0807020",
            INIT_RAM_02 => X"EBF5FAFD7EBF5FAFD7EBF5FAFCFEBF3FAFD7EBF5FAFD7EBF7FBFDFEBF5FBFD7E7F3F9FC6",
            INIT_RAM_03 => X"69B49C6AA550E1245171DD71D96DB6DBAFD7F3F9FDFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_04 => X"140604030180E0604824100803838944805128900A24828940C24838A4924AA5538DE6F3",
            INIT_RAM_05 => X"EBF7FAFD7E7F3F9DC6E36DB6DB6DF6FB7DC6E3F1B8DC6E36DB4DA6CF63B0B75B2D3268E3",
            INIT_RAM_06 => X"EBF5FBFD7EBF7FAFD7EBF5FAFD7EBF3FAFD7EBF5FAFD7E7F5FAFD7EBF5FAFD7EBF5FBFDF",
            INIT_RAM_07 => X"449C564C26534E590381BADE6D369AA9547944DB70B96DB6DBAFDFF3F9FCFF7FBFDFEFF7",
            INIT_RAM_08 => X"C2E16DB65A6D123851100A060481806080401C184C261241C4C2482C9209051389C4A292",
            INIT_RAM_09 => X"EBF5FAFD7EBF5FAFD7EBF5FAFCFE7F1B8DB6DF6DB6DB6DB6DB8DC7E7F3B8DCEDB69B3D96",
            INIT_RAM_0A => X"F3F9FEFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7EBF7FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_0B => X"28920A06134AC8E2AA59289D6EB79B4E592C96491C70379B4DA6AA595B6EB8ED373FAFDF",
            INIT_RAM_0C => X"E3F1B8DB6D767B2D8DC2DB6CB55A24D1E6400C06060301C100A04020144A25130944E261",
            INIT_RAM_0D => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5F9FD7EBF5FAFCFE771B8DB6DB6DB6DB6E371B8FCF",
            INIT_RAM_0E => X"71B8EEB85DB71FAFDFF3FBFDFF7FBFDFEFF7EBF5FAFD7EBF5F9FD7EBF5FAFD7EBF3FAFD7",
            INIT_RAM_0F => X"20120A250309C4C271289C4E27144AA984C279BADF6D289BCE8954AA492492489B4E0703",
            INIT_RAM_10 => X"E371B6DB6DB71B8FCFE36DB4D96CAE170B75B2DB6AB55A24D1A6200C060402818120A251",
            INIT_RAM_11 => X"EBF5F9FD7E7F5FAFD7EBF5FAFD7EBF5FAFCFEBF9FAFD7EBF3F9FD7E7F5FAFC7E771B8DC6",
            INIT_RAM_12 => X"9A44E5913924D2691496452CB85DB71FAFD7F3F9FCFF7FBFDFEFF7EBF7FAFD7EBF5FAFD7",
            INIT_RAM_13 => X"1006030201C100A0401C1A4D25134184D271289C5547169289651389C0E06D289C92CB44",
            INIT_RAM_14 => X"E371F9FCFE771B8DB6DB6DB6DC6E371B8DB6D367B3D85BEDD6EB6DB2D96AB4DA24B16428",
            INIT_RAM_15 => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF3F8DBEDB69B6D9E",
            INIT_RAM_16 => X"89C4DF7349A5128924924928924924B2692C964B2CB96DB71FAFDFF3F9FCFF7FBFDFEFF7",
            INIT_RAM_17 => X"AAD96A944A24B124200C080501810100A061309010289389C4C261449C5A4926930A0703",
            INIT_RAM_18 => X"D36570B75BADF6CB54B25F71BAED76DB8DB6DB6DB6DB6DB6DB4D8EC2DF6DB65B6DB6DB65",
            INIT_RAM_19 => X"EFF9FCFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF1B4DA6",
            INIT_RAM_1A => X"5924944C259349E7249A48DE7039A5524923A25126924AA556892C8A512DB8EDB71FAFD7",
            INIT_RAM_1B => X"B6D96CB5CAA596CB54AA552A9449A49080000C1006051349848061449C4D26148A4512B2",
            INIT_RAM_1C => X"EBF5FAFD7E365B5DAECAE7B0B7DB6DB6994489CEEC95CB2DF72B9ED769B4DA6D367AFB6D",
            INIT_RAM_1D => X"A6D96CB96DB71FAFD7F3FBFDFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7EBF5F9FD7E7F5FAFD7",
            INIT_RAM_1E => X"48AC9547155289A4B2612C994E36138DE724A244DA503925524934A249289449A4B26914",
            INIT_RAM_1F => X"C2DF73B9ECB616CB65A2552A944A25528954AA55289349A44C40180C0E0A051389C4C271",
            INIT_RAM_20 => X"EBF5FAFD7EBF3F9FD7EBF5FAFD7DB69B2DA6BEE36A954AE4F2573BA1D327764A6592A954",
            INIT_RAM_21 => X"A2492691371CD2AB65B6DD6EBB6DB71F9FD7F3F9FEFF7FBFDFEFF7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_22 => X"100A06040492452471512A922895530954D271BCD950B6938E49249A4D1D703924924924",
            INIT_RAM_23 => X"A1D0E994391CAEC923B2592C9A5A2389E6EA79DB6EB449A49249249E492692489B8C3018",
            INIT_RAM_24 => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7E7F5F9FC7EBF5FAFD7DB65B1D96D769A598DBEDB68943",
            INIT_RAM_25 => X"9E4920703AA4D2693C92492593496596AB75B2D96DBA6DB71F9FDFF3F9FDFF7FBFDFEFF7",
            INIT_RAM_26 => X"89C2E172471AA8400018080604824184E27138A4554B2592C954CA79B89D6E36140DE724",
            INIT_RAM_27 => X"D75F6FB6DCF552892B95C8E572395C2A254391C8E4743A65F6592B95BA9C56DB6D522713",
            INIT_RAM_28 => X"F3F9FEFF7FBFDFEFF7EBF5FAFD7EBF5FAFCFEBF3FAFCFEBF5FAFD7EBF5FAFD7E369B0B9E",
            INIT_RAM_29 => X"75C4E0724652C9E70B924921723AA44EA93489DB68944BADB6AB65B2D96EBA6DB73F9FDF",
            INIT_RAM_2A => X"C2DF6996DBED524924A242E071369308B21810080805028944C26138A44E2A25924564D2",
            INIT_RAM_2B => X"EBF5FAFD7E369ADB65B2E9B2B65CB572772B95D92772B95C8E15128540A473BB6E36C964",
            INIT_RAM_2C => X"B6DF71DA6DB73FAFDFF3FBFCFF7FBFDFEFF7EBF5FAFCFEBF5FAFCFEBF5F9FD7E7F3FAFD7",
            INIT_RAM_2D => X"5530922A2593CDA4E36934A27036138E2723A24D249349A4D2A944AA596A94CB6D56AB75",
            INIT_RAM_2E => X"91C8E474495D0E24EAB25B6DB85C2DF6EB75B2D12CB5481AA91240389C51289309410291",
            INIT_RAM_2F => X"E7F3F9FD7EBF3FAFD7EBF5FAFD7E369ADB5CAE6374D6DC2DF677449DD727723A1CAE14E1",
            INIT_RAM_30 => X"B2D528965C2DD6DB85B6DD6DBB6E371FAFD7F3F9FEFF7FBFDFEFF7EBF5FAFD7EBF3FAFD7",
            INIT_RAM_31 => X"75B4922C2592A902B26932964D26144E16E361491E6D261309950392492273485D12B954",
            INIT_RAM_32 => X"A2636474C7548E5743AA3C9D4F291AA5B2E97CD92A965B6D96FB65BEDB6EB85B2CD216C2",
            INIT_RAM_33 => X"EBF5FAFCFEBF3F9FD7EBF5F9FD7E7F1FAFD7E7F5F9FD7EBEDB4D5CB6D531B7DC2DB6C964",
            INIT_RAM_34 => X"71C2E69349E552A944AA492A985BAE16DB136140F0BB6DB71FAFDFF3FBFCFF7FBFDFEFF7",
            INIT_RAM_35 => X"BEDF6EB75BEDF6DB5C9A4D226FB6138994E348ACA06D25144E470B85C9206E371B8DD703",
            INIT_RAM_36 => X"B6CD32D7DBED52893BAE4D34B7D8148E1564CEBA982D185C8D50A8603462702A64D26944",
            INIT_RAM_37 => X"F3F9FCFF7FBFDFEFF7E7F5F9FD7EBF5F8FD7E7F5F9FD7EBF1FAFC7EBF3FAFD7E7F1F6D7D",
            INIT_RAM_38 => X"91BAE171379C0DC6EB654D22734AA512B95492552EB75BEDB6FB4491C931BB6E371FAFD7",
            INIT_RAM_39 => X"58A21948844C0E8954BEE36EB6DC6DF6FB75B2D72271389BCDC71371BCD84D271C4E270B",
            INIT_RAM_3A => X"EBF5F9FCFEBF5F4D96BED533D85B6D528954BEC931B4491BC9C544D2C29C2F2794EDC502",
            INIT_RAM_3B => X"BEE5B1DA6E3F1F9FD7F3F9FEFF7FBFDFEFF7E7F5FAFCFE3F5F9FD7EBF1FAFC7EBF1FAFC7",
            INIT_RAM_3C => X"9A4D226E2613EDA50375B8E49037138DE6D26944E4713AA512893CAA5D6EB85BAE16FB65",
            INIT_RAM_3D => X"B6C8DD564713CECB6475305827044CD2A96DBADB6FB6DC6E36DB6DB2D7249349A4F248EB",
            INIT_RAM_3E => X"EBF3FAFD7EBF1FAFCFEBF5FAFD7EBF5F8FA6CF5B6DB85B6D96895CB6D56DB23A240B4B7D",
            INIT_RAM_3F => X"B2DD70B85C2E172D8ECB6372DB6E3F1F9FD7F3F9FEFF7FBFDFEFF7EBF1FAFD7EBF5FAFD7"
        )
        port map (
            DO => promx9_inst_10_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_5,
            RESET => reset,
            AD => promx9_inst_10_AD_i
        );

    promx9_inst_11: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"AA552A95489C8EB924924D2A9139A38E071391BEE26EB693ADF70375C4E27249A532A93C",
            INIT_RAM_01 => X"CF6BAB94491C8D9544AA48D632BA248EFB5CB2C0D508975596CB75C6E372B8DC6DD6CB6D",
            INIT_RAM_02 => X"E3F3FAFC7E3F1F8FC7E3F1F8FC7E3F1F8FC7E3F1F8FCFE7F1F8FB6A65D68975AADF6697D",
            INIT_RAM_03 => X"75C4E793C9E5527954A25D70B96CB67B3D8ECAE372DA6E373FAFD7F3FBFCFF7FBFDFEFF7",
            INIT_RAM_04 => X"CADB6FB8DC6DB6A93CBADB6CB549A40EA954A25B6A93492492691391B4984EB6538DF713",
            INIT_RAM_05 => X"CF67A9944B6E773B9DBEDF73B03B2552DB54C2CEE052BA25B6CB5CB6D521703AA5B6CB75",
            INIT_RAM_06 => X"F3F9FEFF7FBFDFEFF7E3F1B8FC7E3F1F8FC7E371F8FC7E3F1F8FC6E371F8DC6E7F5FAFCF",
            INIT_RAM_07 => X"9A38DA5546538E271381B8E69249A5329965B2DF70B96CB65B1D85C2E172DB6E371FAFDF",
            INIT_RAM_08 => X"B6D96CB34A25B6FB85CADD6FB6DAE5F6CB6DBEE36895492329E73CA25D6A965A2492A924",
            INIT_RAM_09 => X"E371B8DC6E7F5FAFC7E365B1B149A5D72B44C6DB73B3491B8AB96DCEC8E474491D133B7D",
            INIT_RAM_0A => X"BEDB72DA6DB71FAFDFF3F9FEFF7FBFDFEFF7E371B8DC6E371B8FC6E371B6DC6E371B8DC6",
            INIT_RAM_0B => X"B6D969965AA59669249234A46E37140E072371C4E073491C928944BAE5B2D96CF5F6895C",
            INIT_RAM_0C => X"CED528965925B6FB65B2DB6B96DB6DB6DB6DC6E36DB75BEDB6EB6DB6DF6DAF3592CAA975",
            INIT_RAM_0D => X"E371B6DC6E36DB8DB6E36DB8DC7E7F5FBFCFDB6DAEB85B2DD70B4CBED72896D9DC0E4744",
            INIT_RAM_0E => X"BAE3B3DA6CF5B5D72C713AF4DB6E373FAFDFF3F9FEFF7FBFDFEFF7E371B8DC6E371B6DC6",
            INIT_RAM_0F => X"AA49226AA654D2DB75C2DD6DB44B2DF6EB7581C92891379CD268E3594D216E391CD2893C",
            INIT_RAM_10 => X"C2DB6A96D91C8E4744C6D72FB659A596FB65B2D966965B2DB71B65C2E370B75BEDD6DB7D",
            INIT_RAM_11 => X"E371B8FC6E371B8FC6E371B8DC6E371B8DC6E371B8DCFEBF5FBFCFE3EDB1D85AA616692C",
            INIT_RAM_12 => X"653EE06FB81CD2A934C2E5B2B8ECF67B1B85CB6172DA6E3F1FAFDFF3FBFCFF7FBFDFEFF7",
            INIT_RAM_13 => X"C2E5B2D7DBED1246E3753CE16B279CD2EB9DC75F69913B2DB70B65AA49269349E40D94E3",
            INIT_RAM_14 => X"E36DB2D75C2D96EB9EB6D127754A25B669549A572CB5CAE512DB6DC2DB72D6DBAE174D6D",
            INIT_RAM_15 => X"F3F9FEFF7FBFDFEFF7E3F1F8FC7E3F1F8FC7E3F1B8FC6E3F1B8FC6E3F1F8FD7EFF5FAFCF",
            INIT_RAM_16 => X"B6D9648F3924B1C73489D131B1389BAE4954CF6173DA6D3636DB65B2E174DB6E371FAFDF",
            INIT_RAM_17 => X"B2D96EB75C6E571B9ECB65B0B859A3CD84AA71B2A4754925B6FB9EB6DF6592BAA656EB7D",
            INIT_RAM_18 => X"E3F1F9FD7EBF5FAFCFDB6DB1D759265ADB65CF636A954AE512697DAA552DB6DBADF6DB6D",
            INIT_RAM_19 => X"384932DB6DB73FAFD7F3FBFEFF7FBFDFEFF7EBF5FAFD7EBF5F8FD7E3F1F8FC7E3F1F8FC7",
            INIT_RAM_1A => X"BECB1E70BB6E370B85B6D96495481D52B8FBAE3CE2703AA42E4934B6E373DA6CB61698C2",
            INIT_RAM_1B => X"C2DB6AB7DB6DF6FB7DBADD6DB8DB6E172B85C2E9B2D7DAA34984C25930ACB7DC6E3B2B8E",
            INIT_RAM_1C => X"EBF1F9FCFE7F3F9FD7E3F3FAFDFF3F5F8FC6DB6DB4D85B2CB30B85A25D6996DAE5B6896D",
            INIT_RAM_1D => X"D769B2D9ECF616CB137538F3DB6DB71FAFDFF3F9FEFF7FBFDFEFF7EBF5F9FCFEBF5FAFC7",
            INIT_RAM_1E => X"9A5D74D95CAE3B1D85B6D719564C2E9B2D85C2DB68934A24D2492385C8E17249E4D2176D",
            INIT_RAM_1F => X"BAD56CB55B6D52DB75D35D6CB6DB2E370B75CADD70B85C2E5B0B85CAE170B8589B09C513",
            INIT_RAM_20 => X"E7F5F8FD7EBF5F8FD7EBF5F9FD7EBF5F9FD7E3F3FAFE7EBF5F9DC6DB6DB3D85C2DD6EB6D",
            INIT_RAM_21 => X"85D1227239A4D20713BAE7B0B85CB6372D95C2E3B2DB6DB71FAFDFF3F9FEFF7FBFDFEFF7",
            INIT_RAM_22 => X"C6E5B0B859A2CA477DC2E371B8DC6E373D75B6C8E276DC6E5B2B85CADF70B6DB6D966934",
            INIT_RAM_23 => X"DB69B4DA6CB63AAB85B6CB2CB65BED32CB85C2E36EB54BADF6DB75B6D572B65C2DD70B8D",
            INIT_RAM_24 => X"F3F9FEFF7FBFDFEFF7EBF1F9FC7E3F1F8FC7E3F1B8FC6E3F1F8FC7E3F3FBFD7E7F3B9DC6",
            INIT_RAM_25 => X"BEE370B54A65968913A24D2893C9A4F24944B2EBB3D65C2E3B0B8EC6DB74DB6E371FAFD7",
            INIT_RAM_26 => X"BAE36EB6DBADB73D75C2E170B7D79A8A698DCB67B3D6DC2DB6FB9ECEB2A9954C2E372D9E",
            INIT_RAM_27 => X"E373FBFCFE7F1F8DC6D36DB6D9ED365AEB55C2C52592CB6DD6DB85BEE16997DB6DD6DB9D",
            INIT_RAM_28 => X"CB6174DB6DB71FAFD7F3FBFCFF7FBFDFEFF7E773F8FCFE371B9FC6E371B8DC6E371B8DCF",
            INIT_RAM_29 => X"B2C922765C2E371B85C2DF6EB85C2D9669139248E696DAA4D26913AADB70B85BADF72D96",
            INIT_RAM_2A => X"BADB6DB7DC2DD6EB6DBED56EB6DC2DD70B8DCB65AEB8D75C0ECB96CF6BB3D95B6DF6B975",
            INIT_RAM_2B => X"E36DB7DB6DB6FB8DB6E375F9FCFE371B8DB6DB71B6D9ED365B0B55A26BB0B6DB2DF6EB75",
            INIT_RAM_2C => X"9A6172D6DC2D52CB9ECEE174DA6E3F1F9FD7F3F9FEFF7FBFDFEFF7E371B8DC6DF71B6DBE",
            INIT_RAM_2D => X"CF67B4D8DBED92DB85B2D326965BEDF73D9EAE5972BAECAD1248D2924F2492481C4E7934",
            INIT_RAM_2E => X"71C0F0B75B2E170B75B2DB70B85C2E16DB54BAE16EB7DCAE16EB96CB65B0B7591D12FB95",
            INIT_RAM_2F => X"DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB73F9FCEE3F3B6DC6E36DB8DA6D3616EB44",
            INIT_RAM_30 => X"81C924913B6C4E1723AA4D2EB85BAD9606AA81D973DB6E3F1FAFDFF3FBFEFF7FBFDFEFF7",
            INIT_RAM_31 => X"C6E5B2D659A5F6FBAECF6572BA6C2D12C96DB6D131B6DBAE372B85C2D96DB95C2D968965",
            INIT_RAM_32 => X"E371B6DA6C75D6AAD361245E744BAE16EB85B2E16DB85C2E56FB65B2DD6CB75C6D96DB85",
            INIT_RAM_33 => X"F3F9FEFF7FBFDFEFF7DB6DB6DB6D36DB5DA6DB69B4DA6D369B6DB6E373F8FC6E771B8DCE",
            INIT_RAM_34 => X"BADD72B7DB6DB6A94471D51D7039644E2703B2CD26985BED96A8CA75C0F4DB6DB71FAFDF",
            INIT_RAM_35 => X"B6E16DB6DBECD2A985C7616DB1375B099544CF67B3D9EC2D92C97DB6C4E994CB2D972B7D",
            INIT_RAM_36 => X"E371F8DC6E371B9DCEE36DB4DA6BAD31A6B271B8DA554B2DF6EB85B2DD68985C2E56DB85",
            INIT_RAM_37 => X"81B8F6DB6DB71FAFDFF3F9FEFF7FBFDFEFF7DB6DB6DB6DB6DB5DAED76DB4DAEDB6DB4DB6",
            INIT_RAM_38 => X"B6CB25965BED130B8DBAD96EB65B6DF6DB24B2C8D94AAA64D24934AA512696DC2DD6FB54",
            INIT_RAM_39 => X"BAE370B6DB2E16CB75C2E16AB6D9E40EDB95C2D9584403C9E5124844CD31B96D35B6C94C",
            INIT_RAM_3A => X"DB6DB5DB6DB6DB6DBEE771B8DC6E373F9FCEE36DB4D6DAAD95E703613CEA944B6DD6697D",
            INIT_RAM_3B => X"AA596CB65BADD70B75B6D976DB6E373FAFDFF3F9FEFF7FBFDFEFF7DB6DB6DB6D36DB4DB6",
            INIT_RAM_3C => X"61102077DB6D32994CA244EC96DBEE573D8DBAE9ACB64BED96CB54694D134AA75C0E690B",
            INIT_RAM_3D => X"79D520754B2D12DB6DCADB6DB85BAD96896DB6D96DB65AA4932B96C29408081713CDD4F3",
            INIT_RAM_3E => X"DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DC6E3F1B7DB6E371F9DC6E36DB3D85AAC0DE6B2",
            INIT_RAM_3F => X"B2B4AB8E371BCE7954AE5968954B6D12EB85BEE174DA6E3F3FAFDFF3F9FEFF7FBFDFEFF7"
        )
        port map (
            DO => promx9_inst_11_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_7,
            RESET => reset,
            AD => promx9_inst_11_AD_i
        );

    promx9_inst_12: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"9A1A10292B6D742092612A8914CB6DB65964965328965B6DD72D9EBEDF6DB7DCAD56A924",
            INIT_RAM_01 => X"DB6DB1D96A64B1E6E355492CB65AAE170B65AAE56DB85B2D96CB559A596CB659A40F1D75",
            INIT_RAM_02 => X"F3F9FEFF7FBFDFEFF7DB6DB6DB6DB6DB6DAEDB6BB6DB6DB6DB6DC6E371B7DC6E7F1F8FC6",
            INIT_RAM_03 => X"CF616EB95BEDB689246955226D25544E49449A512A96DAA596CB6DBED972DB6E373F9FDF",
            INIT_RAM_04 => X"BEDB6EB6D9A5B6FB8D38880D20000000003024B28E2CAC6DF6996DB25B6DB54B2E372B95",
            INIT_RAM_05 => X"E3EFB6DC7E3F1F8DC6DB69B2D759A45226EB5940E272489D12896DAA6170B65C2E16DB85",
            INIT_RAM_06 => X"AE5972DA6E3F3FAFDFF3F9FEFF7FBFDFEFF7DB6BB6DB6D76DB5DB6D76BB5DAED76DB6DC6",
            INIT_RAM_07 => X"95E16DB6DAA69B1D85B6E56CB7DC6D96696D81C4EDB2491C2DF6EA89D126954AA552A965",
            INIT_RAM_08 => X"AA5B70B75BAD56CB55A6616DB85B6D52CB8D348C0D2000000000300832912A1B6D52874C",
            INIT_RAM_09 => X"D76BB4DAED76BB6DC6E371B6DDFEBF3F6DB6D365AEB5581CD2B8D26530A06E39A4D2CB24",
            INIT_RAM_0A => X"89D12CB75B2D96AB54AA512EBA6E3F3FAFDFF3F9FEFF7FBFDFEFF7D369B4DAED36BB5DA6",
            INIT_RAM_0B => X"183292481B6DB6C91396512CB3CB6E773D9ECF6172B95BAD971B2381BADD6FB71AC9A4FB",
            INIT_RAM_0C => X"96511C75475BAD13547DDB6897596492AB65AADB72D8EC2DB71B75180C12200000000008",
            INIT_RAM_0D => X"D76BB5DAED36BB4DAED76BB5DAED76DB6DC6E3EFB9FDFE7F1B4D9ECB616DB55AA42D5503",
            INIT_RAM_0E => X"85CF2890B79AA912A271C4EA96DB6D96A965B2D536DA6E3F3FAFDFF3FBFEFF7FBFDFEFF7",
            INIT_RAM_0F => X"2006154B29A8200079693CC6081AA5D5C52BB25B6996D9267B1BA6CF67B2BA6B2DB6A934",
            INIT_RAM_10 => X"B6D56894479DB626F39A4D227346540E88C2594D22723AA44E4924B2D12EB8EC2E572BA6",
            INIT_RAM_11 => X"F3FBFEFF7FBFDFEFF7D769B5DAED76BB5DA6D769B4DAED76DB6DCFE7F1FAFDFE7EDB4D75",
            INIT_RAM_12 => X"B2E7B3D96C2E56CB349A48E07137138D44AA5940EA965B6DB6EB4CAACD2CBA6E3F3FAFDF",
            INIT_RAM_13 => X"89C0E5944BAE16EB855114080B2B6CB1C7036918430B2B6D92576DB2E16CB6D48EBAEB95",
            INIT_RAM_14 => X"EBF5FBFDFE769B1D75AA512495C79C8E068971AC9D765B6C91E75489BCD84A1924D1D734",
            INIT_RAM_15 => X"B2D532BB6E3F3FAFDFF3F9FEFF7FBFDFEFF7D76BB5DAED76DB5DB6D36DB5DAEDB6DB6DC7",
            INIT_RAM_16 => X"B6D92991381E9B1B9DCF69B2B96CF5D6CB549A492A924AA511A4AA6940EA965B6DF6AB65",
            INIT_RAM_17 => X"71A69D75481C0E697575B4DA52481E171D6DC69A00030552A964AA2C800D13CC6C2E876D",
            INIT_RAM_18 => X"D76BB6DB6DB6DB7DC7EBF5FCFD7E369B0B65A24D206CA653ADC7447DB0ACB4481CD2EB75",
            INIT_RAM_19 => X"6132A6965AA596EB65BAD531BC6E3F3FAFDFF3FBFEFF7FBFDFEFF7D769B6DAED769B5DAE",
            INIT_RAM_1A => X"248C1D78DD3532C9759632985546569AEB3CCAE5B4D9EC6DD6CB44B2C4E473C9A4D268FB",
            INIT_RAM_1B => X"44C92A913BACD2896D9E284D2E3692C9E775A240D84CA81C930B96C6D948038000201008",
            INIT_RAM_1C => X"D76BB6DA6D76BB5DAED76DB6DB6DB6DB6DD7EBF9FCFD7E3E5AFB55A244DC713692C902CA",
            INIT_RAM_1D => X"A24D279449A4F2894471C922754B2DD6CB6DBED96FBB6E3F5FAFDFF3F9FEFF7FBFDFEFF7",
            INIT_RAM_1E => X"D365AA8EB3410020000040EC97CBE5930B4C814AD434CAA676898DD367B3D9ECF656CB65",
            INIT_RAM_1F => X"9E4D22713593ADC6D26934A076DC6D55E785C2CD30B65AA5B62744CF63B1B55AA5B6CB9E",
            INIT_RAM_20 => X"F3F9FEFF7FBFDFEFF7DB69B6DAED76BB4DB6D76BB6DB6DB6FB7DCFEBF9FCFD7E3E9ADB55",
            INIT_RAM_21 => X"C2E3B2B85C765B0B65B2DB6A95CAA5527924614922724B2DF70B6DBADD72DB6E3F3FAFDF",
            INIT_RAM_22 => X"B6E16EB96D76172DA6D369B2D9EAE42D424050AA9C52B95D0E24DA89532DB03AE6BA27A6",
            INIT_RAM_23 => X"EBF7FCFDFE3E9B0B65AA4D2270369205656DAA552A92371A0626A279DD648D26542D85AE",
            INIT_RAM_24 => X"BADF6EBB6E3F3FAFE7F7FBFEFF7FBFDFEFF7D76BB5DAED36DB5DB6D36BB6DAEDB6DB6DD7",
            INIT_RAM_25 => X"A65F70B7DD767B1BBECB67B0B9EC2E571D75B6D96CB65B2D528923693099523B2DD6FB75",
            INIT_RAM_26 => X"555969955B29C6074489E16AB75C2D572D95C2E9B4DA6CB676693B712A8C2A171AA55312",
            INIT_RAM_27 => X"D76BB5DB6DB6DB7DCFEBF9FCFDFE7E9B2B6DAA4D2070B81B49E6A16144E07139A451E754",
            INIT_RAM_28 => X"79CD1D723AE5D6EB8DBEDB71DB6E3F1FAFDFF3FDFEFF7FBFDFEFF7D76BB6DA6D76BB4DB6",
            INIT_RAM_29 => X"A6511850261329C52BA65930B95D76371B9EB6E171B6DBAE173D85B2D96CB65B2D128913",
            INIT_RAM_2A => X"9A44D94E385CD268C2B6BCE278DA6491850385DF6A975CF656AB7DC6DF6CB6DC2E9B1B65",
            INIT_RAM_2B => X"D76BB5DAEDB69B5DAED76BB6DB6DB6DB6DC7EBF9FCFE7EBEDB2D85B2D1226FB693CDC6CA",
            INIT_RAM_2C => X"BAD96CB54AA512270389C8E7954B2DB70B75B6E16EBA6E3F1FAFDFF7F9FEFF7FBFDFEFF7",
            INIT_RAM_2D => X"BEE56896DC6E573B8DC6E570B4C752C934E285C2EFBA6D367B3DA6C2D96FB54BAE171D85",
            INIT_RAM_2E => X"B6D96A9037DAC942A271D12B8CA61492EB446142EA934AA5D554AA925925985CF616AB75",
            INIT_RAM_2F => X"F3FDFEFF7FBFDFEFF7D76DB5DA6DB6BB5DB6D769B5DAEDB6DB7DC6EBF7FCFE7EBF1B4D96",
            INIT_RAM_30 => X"CEDB66954BAE171D8DBAD56CB54AA4D248EB693EEA96DBADD70B6DA6D52CBB6E3F3FAFDF",
            INIT_RAM_31 => X"615B68913A6552DB54B2D96EB54B2DB6FB8DC75F70B4C5538A04E2711A1D575CB67B3D85",
            INIT_RAM_32 => X"E7F7FCFE7EFF1F7DA6C2DF69B1371BCD64E365225C4F39A4D102A285C0D84FBB2CF15489",
            INIT_RAM_33 => X"B2D96CBA6DB73FAFDFF7F9FEFF7FBFDFEFF7D76BB5DAEDB69B5DAED76BB5DAEDB6DB6DB6",
            INIT_RAM_34 => X"711A460CAB6E5A897DBED96695CBEDB70B85C2DB6EB75A6D1228F39A5528965B6DD70B75",
            INIT_RAM_35 => X"71A4584C244B48A0916910112AA85CB29965B6D96A96DBEDD6DB8DC2E370B6495C2DE4EA",
            INIT_RAM_36 => X"D76BB5DA6D76DB6DB6E375FAFE7EBF3F8DB6CB6170B4485B4942D289B8DC6896949288E3",
            INIT_RAM_37 => X"89D52CB6DBADD6EB6DB6DB6DBA6E373FAFDFF3FDFEFF7FBFDFEFF7D76BB5DAED76BB5DAE",
            INIT_RAM_38 => X"C6DF6FB64A64AE992C81920308981DB6CB6DAE5124765B2E173D8DB6D96CB4DAA4D22724",
            INIT_RAM_39 => X"5540EB8D2BEB4A88B281A25128948A44D26971A0554E279D3258CA79D31E734B6D12DB7D",
            INIT_RAM_3A => X"D76BB5DAED76BB5DAED76BB5DAED76BB5DB6E375FAFE7EBF5F9DB6D369B0B4D89BCDA4B2",
            INIT_RAM_3B => X"BAD36A9249240DE6A29E596EB75BEDB6EB65AA5570BB6DB71FAFE7F7FDFEFF7FBFDFEFF7",
            INIT_RAM_3C => X"924D2DB85B25B6DB6DC2D92996CA1D32574C5510090202040E472395C8E896DC2E172B85",
            INIT_RAM_3D => X"DB6DB2D7589C0D64F3924B26995B2D12CB34B2D11E72C926370B4DB6BAE07859E5B6794C",
            INIT_RAM_3E => X"F3FDFEFF7FBFDFEFF7D36BB4DA6D369B4DAED769B5DAEDB6BB5DB6DB75FBFE7F3F5FBFCF",
            INIT_RAM_3F => X"38B8A5985B6E571D8EB6D5248E375C4E6944A2596CB75C2E16DB6DAAD130BB6DB73FAFE7"
        )
        port map (
            DO => promx9_inst_12_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_9,
            RESET => reset,
            AD => promx9_inst_12_AD_i
        );

    promx9_inst_13: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"6542E0765BAD970B34C2DB65965B6D52CB6DB6DB6F943A1D0E991265140D089280A154D3",
            INIT_RAM_01 => X"DB71FAFE7EFF9FAFCFE3F1B6D8EA6B4E071392552298DAADD6AB2CC2E16CB4489ACA0689",
            INIT_RAM_02 => X"B2D570BB6E3F1FAFE7F7F9FEFF7FBFDFEFF7D369B4DAED369B5DA6D36BB5DAED76BB6DB6",
            INIT_RAM_03 => X"859A0E040180A0606840C0EC94CBEE5B1D85B2CF2270375C4EA96DB2D96A965B2D96DB75",
            INIT_RAM_04 => X"B2E1688F35140E6954B2D969B6DB6DB6CB7DBED96DB659A5B6FB8DBAD96DB43A1D329913",
            INIT_RAM_05 => X"D369B5DAED76BB5DA6DB71BAFD7EBF9FBFD7E7F3F8DA6AAB8B2D34AAC4E690BAA536AB75",
            INIT_RAM_06 => X"B6DB6CB65AA5B6CB6DB2CD30BB6E3F1FAFE7F3FDFEFF7FBFDFEFF7D369B4DA6D769B5DA6",
            INIT_RAM_07 => X"B6D52A9238144E0703611A11271243CE47236144EC97DC2E7B3D85AA511C6D289CD2A965",
            INIT_RAM_08 => X"712859524695F6890B8A246274CAA5530B85C2E3B2D75CADB6EB55B6D56FB85B6E570B75",
            INIT_RAM_09 => X"D369B4DA6D369B4DAED36BB4DAED76BB6DB6DB6DBAFD7EFF7FBFD7EFF3F8DB6C75D626C2",
            INIT_RAM_0A => X"9A44E26EBAA552CB65B2D96AB549A5129B6DAACB31DB6E3F1FAFE7F3FBFEFF7FBFDFEFF7",
            INIT_RAM_0B => X"C2EFAEB34B6D52A964A64AD94AA7542994EA341C542EAA2572A95C9A4D30B8DCAE5B2D55",
            INIT_RAM_0C => X"EBF5F8DB6C2C516513653AD64D29A3CDA4FB593492450A25369B65B2E570B75BAE5B2D85",
            INIT_RAM_0D => X"F3FDFEFF7FBFDFEFF7D769B4DA6D769B5DA6D36BB4DAED769B5DB6DB6DB8FD7EBF7FBFE7",
            INIT_RAM_0E => X"B2CD2DB9EC6E5ADB2C9A4926944AA552A96DB2D96AB449640E294CA6C0EEBB6E3F3FAFE7",
            INIT_RAM_0F => X"4938E6934BAE172D96D7616B93C91B4994814492112AA61329C4C244AAA776DBADB6DB6D",
            INIT_RAM_10 => X"DB6DB8DD7EFF7FBFE7EBF5F8FB6C2C5206E37DCD2A934924D1C6C2AA49258EBA2329A6AA",
            INIT_RAM_11 => X"8A3CF0BB6E7F3FAFE7F3FDFEFF7FBFDFEFF7D36BB5DA6D769B5DA6D76BB4DA6D76BB6DB6",
            INIT_RAM_12 => X"B25F70B96CF6370B85BAD96FB96CF656CB2C9A44E6965B2D52DB65AAD5289138E3CD54E3",
            INIT_RAM_13 => X"B2D52CB4481BAD44C265226A99EC2E573D54719C45020001E5128944C0994A960CAE594C",
            INIT_RAM_14 => X"D76BB5DA6D369B5DA6DB6DB8DD7F3F5FBFDFEBF5F8FB6BAC4E4944B2DF6CB54B6D528944",
            INIT_RAM_15 => X"AA51228F361348E29269B8EDBC7E7F5FBFE7F3FDFEFF7FBFDFEFF7D76BB5DAED76BB5DA6",
            INIT_RAM_16 => X"AE5F6C92B6532A996DC6E7B2D96D365B0B85C2DD70B9EC2CD2592C89C92795CAA596CB54",
            INIT_RAM_17 => X"9A552CB65CAD96AB44B6D9669449A511C7139E532DB85BAE9A884828184E271140007123",
            INIT_RAM_18 => X"D76BB5DAED76BB5DAED76BB4DAED769B5DB6DB6DB6DD7EFF7FAFD7EBF5F8FA68A40E075C",
            INIT_RAM_19 => X"AA512A965B2D96CB549A44D64AA49248A26130A4AEBB6E3F5FBFE7F3FDFEFF7FBFDFEFF7",
            INIT_RAM_1A => X"8E34D12B2591E400B2B2DB68744A638A5703AE5B73D7DD369B2D95C763B3D85AAC925954",
            INIT_RAM_1B => X"E7F3F6D7D79B4944E3AADF6CB85B2D96596DAAD96EB54A24D25955A25B71B75B2BACD0A2",
            INIT_RAM_1C => X"F3FDFEFF7FBFDFEFF7D76FB7DBEDF6FB5DBED76BB4DA6D36BB4DB6DB6DB6DC6EFF7F9FCF",
            INIT_RAM_1D => X"D367B1D85B2D128965BADB6A965B2D5689449A3CD5461281C5247128AAAEBB6E3F5FBFE7",
            INIT_RAM_1E => X"C2D968985B2920A089000000010493ACC2719A676474CB251286AA9A44F0B75D365B5D85",
            INIT_RAM_1F => X"DB6DB6DC6EBF9FAFC7E3E9A890381B8E692CC2E16DB85B6DD6CB54B6D32892CA2552396D",
            INIT_RAM_20 => X"553CEEBB6E3F5FAFE7F3FDFEFF7FBFDFEFF7DF6FB7DBEDF6FB7DAED76BB5DA6D36BB6DB6",
            INIT_RAM_21 => X"89D131B75CF6174DA6CF65AEB65AAD96DB65BADB6DB7DB2D52A9249A309244828A04E291",
            INIT_RAM_22 => X"C2DB68944A25D71B65AA552A975699211200000000000142A9543089E16992C9A5725913",
            INIT_RAM_23 => X"DF6BB5DAED76BB4DB6DB6FB6DC6E3F5FAFCFD3616490389D573D75AAD56CB65B2D56EB65",
            INIT_RAM_24 => X"81B8CC26938A4554D2593CEEBB6E3F5FCFE7F3FDFEFF7FBFDFEFF7DF6FB7DBEDF6FB7DBE",
            INIT_RAM_25 => X"92636574CB6D96FB4C925D6EB75D765B4D9EC6E170B6DB2D56EB75B6DD6EB6DB2CD2A913",
            INIT_RAM_26 => X"92596DB75BADD70B4C9A596AB65AAD970B659A5D6DB44550C13400040000010042455430",
            INIT_RAM_27 => X"DF6FB8DBEE371B8DBEDF6BB5DAED769B6DB6DB6DB6DC6E775FAFCFC2D11C703B2E16597D",
            INIT_RAM_28 => X"BADD6DB65B2D128924692C934AA6138DC6CA653CF1DA6E7F5FBFE7F7FDFEFF7FBFDFEFF7",
            INIT_RAM_29 => X"9A3AC001028AC8D289AE5F6072BA65B6DB75A265B2D65D369B2D96CAE170B85B2DB6CB6D",
            INIT_RAM_2A => X"81C0E8996C765AEB7DC2DB71B6DBEDF6AB4DC2D128975B6D32A944AE5B70B75508811292",
            INIT_RAM_2B => X"F3FDFEFF7FBFDFEFF7E371B8DC6E371B8DC6DF6DB5DAED76BB6DB6DB6DB7DC6E773F8F96",
            INIT_RAM_2C => X"C6E16CB6DB6D96CB6DB2DB6CB55B2D12692471B4944CA65349C6E3654531DB6E3F5FBFE7",
            INIT_RAM_2D => X"B2D96CB6D92140F2CA651E4A2926534C60C2B2D52272CB6DB6DB6D44E5B4D44CF65B3B7D",
            INIT_RAM_2E => X"DB6DB6DC6E373B6D2479D973D96D3596CB7DAE572CB95A25570B34B2D965965B2D56A955",
            INIT_RAM_2F => X"694D32DB6E3F5FBFE7F7FDFEFF7FBFDFEFF7E7F1B9FC6E7F3F8DC6DF6FB5DAED76DB6DB6",
            INIT_RAM_30 => X"89E7B5D44C6E7AFB6DBEE16CB54A6D12AB44A6512994DAACD24913592C934AA6138DC6E3",
            INIT_RAM_31 => X"BAD96396DA6D12CB75B6DB70B75A21A460AA69BCDC6CA611419554A64B2592C81D72FB75",
            INIT_RAM_32 => X"DF6DB7DAED76BB6DB6DB71B8DC6E76DA58F3CAE7ADB85C2DF6DB65AA552CB85C2D36DB55",
            INIT_RAM_33 => X"79C0E26EB79B4984B2655532DB6E3F5FCFE7FBFDFEFF7FBFDFEFF7EFF3F9FCFE7F3F9FCF",
            INIT_RAM_34 => X"81D92996D965971B85C6E7B4D96C6E170B95B2DB6AB55AAC4E592CA24D2CB34A24D20703",
            INIT_RAM_35 => X"AA5B66985CAD52CB6DB6D96996DA25970B55AADD6CB55B6B0994D218164A2593438B5D9E",
            INIT_RAM_36 => X"E7F3F9FCFEFF3F9FC6DF6FB7DAED76FB6DB6DB71B8DC6E7CB24996C2E5B0B85C2D96A98D",
            INIT_RAM_37 => X"964D28954A248DF7249A44DF6F365349C70371CD33DB6E3F5FCFEFF3FDFEFF7FBFDFEFF7",
            INIT_RAM_38 => X"B6CB24965C2E7AEB4CB24B2C97DB6DF71BA6CAE9B5D9EC6DF72D85A25366934963CE0724",
            INIT_RAM_39 => X"B2E7B5D85C2E5ADB54B6CD2A985BAE16CB6DAAD56CB75B6DB6DB75BADB6EB75B6D128944",
            INIT_RAM_3A => X"FBFDFEFF7FBFDFEFF7EFF7FBFDFEFF7FBFCFE36FB7DAEDB6DB6DBEDB71B9FC68A65B2D75",
            INIT_RAM_3B => X"C2CD124E392309A534A24D2694489C8EA9449E492270379BCE07036944F4DB6E375FCFE7",
            INIT_RAM_3C => X"B2D96DB6DA2349E75CBAE3B4D9ECF616B944AE552DB8DB2DB6B96DCF67B5DA6CAE36FB85",
            INIT_RAM_3D => X"E371F8D55CADD74D6DCB67B2D85B2E7AFB6DAA592EB75CF5D6DB65B2D36A96DB2D571B75",
            INIT_RAM_3E => X"71C0F2DB6E375FBFE7FBFDFEFF7FBFDFEFF7EFF7FBFDFEFF7FBFCFE36FB7DB6DB6DB6DB6",
            INIT_RAM_3F => X"CAE572D8EBAE170B75A240D84D369225A5139A59679249E552A954A248E171381C0E06F3"
        )
        port map (
            DO => promx9_inst_13_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_11,
            RESET => reset,
            AD => promx9_inst_13_AD_i
        );

    promx9_inst_14: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"BAD570B75AADD6EB75B6DD6FB5481B0A0765C2E174D96CADF6C964B6D334B7DB2552FB5C",
            INIT_RAM_01 => X"E7EFB7DB6DF6DB7DC6E76FB2B9ECF5970B7DBADD73D55BEE7AB97DB25970B8ECB5F73B55",
            INIT_RAM_02 => X"91C4E271381C0E070379C2F4DB6E3F5FBFE7FBFDFEFF7FBFDFEFF7EFF7FBFDFEFF7FBFCF",
            INIT_RAM_03 => X"B2DB6FB5495D96995CA2616FB6DCB5D6CB2C964D1A4B244A4585039A4F2893CAA596A954",
            INIT_RAM_04 => X"91E775D9DA2572DB6DB2DD6DB2CA2596EB85C2DD6DAEB6932A076DB6E372B8DBADF6FB6D",
            INIT_RAM_05 => X"EFF7FBFDFEFF7FBFDFE36FB7DB6DF6FB6DC6C2E7B3D9EB2E373D8DC2DF74D9EAE636DB6D",
            INIT_RAM_06 => X"924F269249A552A93491CF2691381C0DE70379C4F2DB6E375FCFE7F3FDFEFF7FBFDFEFF7",
            INIT_RAM_07 => X"AAE5B2D6DB6D532B65CF59689139A572A954B2DB6A985A24D26955923AE68AA489852303",
            INIT_RAM_08 => X"D75F6B96DB6DD6898DAE532DB5CA2492B9349A596B94485D52AB8DC2DD6EB4475B8DC724",
            INIT_RAM_09 => X"FBFDFEFF7FBFDFEFF7F3F7FBFDFEFF7FBFDFE7EFB7DBEDF71B6D4CCF69B3D75C2E7B0B9E",
            INIT_RAM_0A => X"71CB184B248A4564E39249269249E5126913AA512691381BCE071389CD32DB6E375FCFE7",
            INIT_RAM_0B => X"BEDF70B6DAA40DD713A2596DB55C2E170B96C2DF6B954BEE36EB6DAE596A965AA44E070B",
            INIT_RAM_0C => X"D36370B95C2E5ADB96CF5F647A6B6E36697DBEE36B954B6C0EA965AE5F66954A25968955",
            INIT_RAM_0D => X"9A5134DC6E377FCFEFFBFDFEFF7FBFDFEFF7EFF7FCFDFEFF7FBFDFE7F1B8DBEDF6BA59A6",
            INIT_RAM_0E => X"92512694479C4E0703AE491A6CA5538D12D3A24D2793CA25128944AA552792C89C4E272C",
            INIT_RAM_0F => X"BEDB6DB6DBAD968975B2DB6FB7DB6DB6DB239A492A94496556DB6DAAE76FB6DA2596CB3C",
            INIT_RAM_10 => X"E7F3F7DBED74735D96C2E7B2D85CF636FBAEBEDB6B97DC6D52B98DBED32C96DAE40EB97D",
            INIT_RAM_11 => X"AA5526934964B269349A5974DB6E7F7FCFE7FBFDFEFF7FBFDFEFF7F3F9FCFE7EFF7FBFDF",
            INIT_RAM_12 => X"89D52CB54B6D5249659244EFB0B92636070389C0DA6E371A89551379C4E2734A2512A954",
            INIT_RAM_13 => X"BEEBB4D9DAE6372D96C2E170B8DCADF6DB65BEDF70B75AAE16AB8DBEDB6DB65AA4B26903",
            INIT_RAM_14 => X"F3F9FCFE7F3F7FBFDFE7F1B7DBEBAE9B3D9ED367B7D96CF67AFB65C6DB6B96DC6DB71B9D",
            INIT_RAM_15 => X"71BCE2754AA5128944A24F269349A4B2692489C4F4DB6EBF9FDFE7F3FDFEFF7FBFDFEFF7",
            INIT_RAM_16 => X"A25526954A25126944A244E8924A2552491389C2E177D81BEE070385D51F713694D184C2",
            INIT_RAM_17 => X"C6E776DB6E373F9DDFE76DB5DA6CF67B3D95CAE7B1D85BAE170B85C2E171B75B6D96AB44",
            INIT_RAM_18 => X"FBFDFEFF7FBFDFEFF7F3F9FCFE7EFF7FBFDFE7EFB7DAECF6BB4D85D36BB3D96BEE573D9D",
            INIT_RAM_19 => X"7DBADE73C7DB0A68B25934A2724A24D26954A251299349A4D27924755B75DC6EBF9FCFF7",
            INIT_RAM_1A => X"BADD6DB75BAD9689549A4B2692C9A4D2A944964928944A24D2692C9A49227249A3ADF6F3",
            INIT_RAM_1B => X"D36BB2D9ECF6BB5DAEDB69B4DB6DB73B9DD7EFF1B6DA6D369B3D9ECB6170B85B6DD6CB65",
            INIT_RAM_1C => X"556174DC6EFF9FCFEFFBFDFEFF7FBFDFEFF7F3F9FCFE7F3F7F9FCFDF6FB5DAECF69B4DAE",
            INIT_RAM_1D => X"A651269449645268EB71BADC6E39A3ADC71361309E713A24D2693CA2512993489CD24713",
            INIT_RAM_1E => X"DF6DB6DAED36BB4DA6D367B0B85BADD6EB7DB6DD6CB54A65728954A25329944A6D12AB55",
            INIT_RAM_1F => X"DF6BB5D9ECF67B3DA6CB65B2DA6CB65B4DA6D369B4D96CB6BB5DBEE3F5F9FC6E36FB7DBE",
            INIT_RAM_20 => X"9E4D2171389C4DE6C271E374DCEEBF9FCFE7FBFDFEFF7FBFDFEFF7F3F9FCFE7F3F5F9FBE",
            INIT_RAM_21 => X"B6DD6EB6DB2D56CB6DBAD568955AA4D2691381B8DC56D613AD84D2612A9E6F39A4D2793C",
            INIT_RAM_22 => X"D371FBFDFEFF9FAFD7EBF5FAFCFEFF3F9DC6DB69B4D96CB67B1D85C76170B75C2E16DB75",
            INIT_RAM_23 => X"F3F9FDFE7F3F5F9FC6DF6BB5DA6D367B3D96CB65B4D96CB69B2D96CB65B2D96CB65B3D9E",
            INIT_RAM_24 => X"71B4A68E39A4B2693C924D2590381BCE270389E574DC7EBFBFCFE7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_25 => X"D365B2D96C765B2D96C763B0B85BADD6EB6DBED96CB54BAD56896DA249216E3A234A16C2",
            INIT_RAM_26 => X"DB6BB4DA6D369B4DA6D36BB8DDFEFF9FCFE7F3F7FCFDFEFF7F9FC7E76DB6DB6D36BB4DA6",
            INIT_RAM_27 => X"FBFDFEFF7FBFDFEFF7F7F9FCFE7F3F5FBFDFDF6FB7DBED76BB5DAED76BB5DAEDB6DB6DA6",
            INIT_RAM_28 => X"AA512491379C2D84D26138D64D29A51289349A4F2691381C0E071389E172DC7EFF9FCFEF",
            INIT_RAM_29 => X"E7F3F9DCEDB6DB6DB6DB6DB6DA6D36BB4DA6D365B3D96C76170B75C2DB6DB6DBAD96CB65",
            INIT_RAM_2A => X"E36DB8DB6E36FB8DC6E371B7DB6DF6FB7DBEDF6FB6DB6E3F5FBFE7F3F9FBFDFEFF7FBFCF",
            INIT_RAM_2B => X"926172DCFEFFBFCFE7FBFDFEFF7FBFDFEFF7F7FBFCFEFF3F5FBFDFE7F3F9FC6E36FB8DC6",
            INIT_RAM_2C => X"C2E16EB75BADD6FB65B2D72893C89C0E78C26134984C2964D26934AA512793481BEE0713",
            INIT_RAM_2D => X"EFF7FCFE7EFF7FAFD7EBF7FAFCFE7F3B9DCEE773B8DC6DB6DB6DB6DB69B4DA6CB67B2D9E",
            INIT_RAM_2E => X"EFF7FBFCFEFF3FAFC7E7F1F8FCFE7F3F9FD7E7F5F9FD7E7F3F8FCFE3F1B8DC6E371F9FD7",
            INIT_RAM_2F => X"A251269247144E4934A25D74DC7EFFBFCFF7FBFDFEFF7FBFDFEFF7F7FBFDFEFF3F9FBFDF",
            INIT_RAM_30 => X"DB6DB6DA6D369B2D85CB65B2D85C2E5AEB75B6E16CB549E48DE713612C9C6D2964D26934",
            INIT_RAM_31 => X"EBF5FAFC7E7F3FAFCFE7F5FAFD7EBF5FAFD7EBF5FAFD7EBF3F9FCFE7F3F8FC7E771B9DC6",
            INIT_RAM_32 => X"F7FBFDFE7F3F9FBFDFEFF7FBFDFEBF3FAFD7EBF5FAFD7EBF5FAFDFEFF7FBFD7EFF7FAFDF",
            INIT_RAM_33 => X"75B0964D28A5128934A255268F381CF2693C925B73DC7EFFBFCFEFFBFDFEFF7FBFDFEFF7",
            INIT_RAM_34 => X"EBF5FAFCFE7F5FBFCFE7F3B8DB6DB6DB6D96D369B4DA6CF63B1B85B6DD70B65AA4F24903",
            INIT_RAM_35 => X"EFF7FBFDFEFF7FBFDFEBF7FAFD7EBF5F9FD7EBF3F9FDFE7F3F9FDFEBF7FBFDFEBF5FBFD7",
            INIT_RAM_36 => X"FBFDFEFF7FBFDFEFF7F7FBFDFEFF7FBFCFDFEFF7FAFD7EBF5FAFD7EBF5FAFD7EFF7FBFDF",
            INIT_RAM_37 => X"C2DF6EB7DB2D52791379B89C6B279C929954AA552690381C8E47349E5974DCFF3FBFEFE7",
            INIT_RAM_38 => X"EFF3F9FDFEBF5FAFDFEBF7FAFD7EFF7FAFDFE7F3F9FCEE371B8DB6DF6FB6DAED367B4D8D",
            INIT_RAM_39 => X"EBF5FAFD7EFF7FBFDFF3F7FBFE7EFF7FCFDFEFF7FAFD7EBF5FAFD7EBF5FAFD7E7F3FBFCF",
            INIT_RAM_3A => X"A25534DCFEFF9FEFE7FBFDFEFF7FBFDFEFF7F7FBFDFEFF7F9FBFDFEFF7FBFD7EBF5FAFD7",
            INIT_RAM_3B => X"E771B6DC6DB69B4DAECB616FB65BED52893485BCDA4C279D128955AA5524924924F2793C",
            INIT_RAM_3C => X"EBF5FAFD7EBF5FAFD7EBF3F9FCFE7F3F9FD7EBF7FAFDFEBF7FAFDFEBF5FBFCFE7F3F8FCE",
            INIT_RAM_3D => X"EFF7FBFD7EBF5FAFD7EBF5FAFD7F3F7FBFDFEFF7FBFDFEFF9FBFDFEBF7FAFD7EBF5FAFD7",
            INIT_RAM_3E => X"AA55289549A4D2493C9A5534DCFEFF9FDFF7FBFDFEFF7FBFDFEFF7F7FBFDFEFF7F9FCFDF",
            INIT_RAM_3F => X"EFF5FAFD7EBF7F9FD7EFF3F9DCEE76DB6DA6D363B0B75B6DB6A93C9240DD6F389D129954"
        )
        port map (
            DO => promx9_inst_14_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_13,
            RESET => reset,
            AD => promx9_inst_14_AD_i
        );

    promx9_inst_15: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"EBF7FAFDFEBF5FAFD7EFF5FAFE7EBF5FAFD7EBF7F9FCFE7F3F9FCEE773F9FCFEBF5FAFD7",
            INIT_RAM_01 => X"F7FBFDFEFF7F9FCFDFEFF7FAFD7EBF5FAFD7EBF5FAFD7EFF5FBFDFEFF5FBFDFEFF7FBFDF",
            INIT_RAM_02 => X"9A42DE6E381CD28954AE572B954AE512A954AA5576DCFF3F9FDFE7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_03 => X"E773B8DB6E371B8DC6E773FAFCFEFF5FAFD7E7F5FAFD7E7F1F8DB6D365B2D85BADB6CB44",
            INIT_RAM_04 => X"EFF7FBFD7EFF5FAFD7EBF5FBFDFEBF5FAFD7EBF5FBFE7EBF5FAFD7E7F5FAFD7E7F5FBFC7",
            INIT_RAM_05 => X"FBFDFEFF7FBFDFEFF7F7FBFDFEFF7FBFCFDFEFF7FBFCFE7F5FBFDFEBF7FAFD7EBF5FAFDF",
            INIT_RAM_06 => X"E371B5D9ECADD6DB54AA44E070389C92AB54A2552CB65B2DB6CB44B2DB74DC7EFF9FEFF7",
            INIT_RAM_07 => X"E3F1FAFD7EBF5FBFCFE7F3B8DC6E371B8DB6DF6DB6DB6DB6DB6DCFE7F5F9FD7EBF3F9FCE",
            INIT_RAM_08 => X"E3F3FAFCFEFF5F9FDFEBF3FAFCFEBF7FAFDFEFF5FBFDFEBF5FAFD7EBF7FAFDFEBF5F9FC7",
            INIT_RAM_09 => X"AAD574DCFF3FBFCFF7FBFDFEFF7FBFDFEFF7F7FBFDFEFF7FBFBFDFEFF7F9FC7E3F3F8FCF",
            INIT_RAM_0A => X"CF69B5DB6E3F1F8FCFE3F3B8DB6D36570B6DAA512270392512B965AA556DB65AA4928965",
            INIT_RAM_0B => X"EBF7FAFE7EBF5FAFC7E371F8FCFE7F5FBFCFEFF3F8DC6E7F1B8DC6E36DB7DBEDB6DB6DA6",
            INIT_RAM_0C => X"EFF7FBFC7E7F3F8FCFE3F3FAFCFE7F5FAFD7EBF5FBFD7E7F3FAFD7EBF5FBFDFEBF5FAFD7",
            INIT_RAM_0D => X"B6D32A9548A349852481C0F4DC7EFF9FCFF7FBFDFEFF7FBFDFEFF7F7FBFDFEFF7FBFCFDF",
            INIT_RAM_0E => X"E36DB6DB6DB6DB6DB6D76BB4DA6CF65B4DB6DB71B8DB6DB69B2D7DB2D1249349A512CB65",
            INIT_RAM_0F => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E3F1F8FC7E3F3FAFCFEBF5F9FCEE373B8DC6",
            INIT_RAM_10 => X"F7FBFDFEFF7F9FCFDFEFF7FBFD7EBF3F9FD7E7F5FAFD7EBF5FAFD7EBF5FAFD7EBF5FBFD7",
            INIT_RAM_11 => X"BAD968924A2556DB65AE51289349230954AA613CF4DCFF3FBFCFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_12 => X"E7F5F9FCFE7F3B9DCEE371B6DB6DB6DB7DBED36BB5DAED36BB3D8DC6E373DB6DB6DB2D96",
            INIT_RAM_13 => X"EBF5FAFDFEFF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF3F9FCFE3F3F9FCF",
            INIT_RAM_14 => X"FBFDFEFF7FBFDFEFF7F7FBFDFEFF7FBFCFDFEFF7FBFD7EBF5FAFD7E7F5FAFD7EBF5FAFD7",
            INIT_RAM_15 => X"CF636FB7DCF69B4DA6CB616CB5496596DB65B2D32894491C0E2703965132DCFF3F9FEFF7",
            INIT_RAM_16 => X"E7F1F8FCFE3F3F8FC7E7F1F9FC7E7F3F9FC6E771B6DC6DB6DB6DB6D76DB6DAED76BB5D9E",
            INIT_RAM_17 => X"EBF3F9FCFE7F5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFCF",
            INIT_RAM_18 => X"A25372DCFF3F9FCFF7FBFDFEFF7FBFDFEFF7F7FBFDFEFF7F9FBFDFEFF7FBFD7EBF5FAFCF",
            INIT_RAM_19 => X"D76BB5DAED369B5DA6CF67B1B7DBAE372D96CF616EB65AAD56DB65B2DB6CB55B2D128944",
            INIT_RAM_1A => X"E7F3F9FC7E3F1F8FC7E371F8FC6E371B9DC6E371B8DC6E371B8FD7E7F3B8DB6E36DB6DB6",
            INIT_RAM_1B => X"EFF7FBFCFEBF3F9FCFE7F3FAFCFE7F3F9FD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E3F1F9FCF",
            INIT_RAM_1C => X"B2DD6FB7DB6D968924A65D71DCFF3F9FEFF7FBFDFEFF7FBFDFEFF7F7FBFDFEFF7FBFCFDF",
            INIT_RAM_1D => X"E3F3F8FC7E771B6DB6DB6BB5DAED76BB5DAED369B3D95C6D96FB95CF63B0B6DAAD56AB65",
            INIT_RAM_1E => X"E7F3F9FCFE7F1B9FC6E7F1B9FC6E7F1B7DC6E36FB8DBEDF6FB7DBEDF6FB6DB6DB6DB6DC6",
            INIT_RAM_1F => X"F7FBFDFE7F3F9FBFDFEFF7F9FCEE7F3B9DC7E773B8FCEE371B8DCFE7F3F9FCFE7F3F9FCF",
            INIT_RAM_20 => X"C2E571B85B2D328965BADD70B6DB6DB6A944AA4D30BCFF3FBFCFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_21 => X"D369B4DA6D369B4DA6DB71B9FCFE7F1F9DB6DF6DB6DAED769B4DAED769B4D9ECF5F6DB85",
            INIT_RAM_22 => X"DF71B8DC6E371B7DBEDF6FB7DBEDF6FB7DBEDF6FB7DB6DF6DB7DAED769B5DAED769B4DAE",
            INIT_RAM_23 => X"FBFDFEFF7FBFDFEFF7F3F9FCFE7F3FBFBFDFE7F3F8DBEDF6FB7DBEDF6FB7DBEDF6FB7DC6",
            INIT_RAM_24 => X"D369B3D9ECF65B2B65BEE172B85BAD966944B6DF6EB4496492A9548E4530BD7F3F9FEFF7",
            INIT_RAM_25 => X"D36BB4DAED369B4DA6D369B4D9ECB67B3D96CF69B9DD7EFF3F8FCEE371B6DAED369B4DAE",
            INIT_RAM_26 => X"D76DB5DAED76DB6DB6DF6FB7DBEDF6FB7DBED76BB5DAED76BB5DAED76BB5DAED36BB4DAE",
            INIT_RAM_27 => X"AADB71DD7F3F9FEFF7FBFDFEFF7FBFDFEFF7EFF5FCFE7F3F7FBFDFE7F1B6DBEDB6BB5DAE",
            INIT_RAM_28 => X"E771B6DBED76BB4DAED369B3D9ECF67B2B75B2E170B95C2DB68944A65B6EB75AAD52CB54",
            INIT_RAM_29 => X"D76BB5DAED36BB5DAED76BB4DA6D369B4DA6CB69B4D9ECF65B4D9ECF67B6DD7EFF5FAFDF",
            INIT_RAM_2A => X"E7F1B7DB6DF6BB5DAED76FB5DAED76BB5DAEDB6FB7DBEDF6BB7DAEDF6BB5DAED76BB5DAE",
            INIT_RAM_2B => X"A2512AB75BEDD6FB85C2E3B2DD7F7F9FCFF7FBFDFEFF7FBFDFEFF7EBF5FAFDFEFF5FBFDF",
            INIT_RAM_2C => X"D369B6DC7EFF5FAFCFE7F3F9DC6DF6FB6DA6D369B4D9ECF67B2D9DBEDF71B8DC7616DB4C",
            INIT_RAM_2D => X"DF6FB7DBEDF6FB7DB6DF6DB7DB6D76FB5DAED76BB5DAED76BB5DA6D369B4DA6D36BB4DA6",
            INIT_RAM_2E => X"EBF3FAFDFEFF7FAFCFE371B7DB6DF6DB7DB6DF6DB6DBEDB6FB7DBEDF6FB8DBEDF6FB7DB6",
            INIT_RAM_2F => X"CADB70B8DC6E16EB659A4D2593496512CB7DC2E3B4DD7F3F9FEFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_30 => X"DF6FB7DBEDF6FB6DB6DB6DB6DC6E775FAFD7EFF5FBFCFE771B7DAED76BB5DA6D367B3D9E",
            INIT_RAM_31 => X"E7F3F9FCFE7F3F9FCFE7F1B9FC6E7F1B9FCFE371B8DBEDF71B7DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_32 => X"FBFDFEFF7FBFDFEFF7EBF5FAFD7EBF5FBFDFEBF3F9FC6E773F8DCFE7F1B9FC6E7F3F8DCF",
            INIT_RAM_33 => X"DB69B4DA6D369B3D9ECF6370B8DC2E3B0B6DA24D24934924920744BAE5B4DD7F3FBFEFF7",
            INIT_RAM_34 => X"E3F1F9FC6E771B9FCFE7F1B9FCFE371B9FC6E371B8DC6E773F9FDFEBF7FAFD7E7F3F9DB6",
            INIT_RAM_35 => X"E7F3FAFCFE7F5FAFDFEFF5FBFDFEFF3F9FCFE7F3FBFCFEFF1FBFC7E7F3FBFC7E7F1F8FCF",
            INIT_RAM_36 => X"BAE5B6DDFF7F9FEFF7FBFDFEFF7FBFDFEFF7EBF5FAFD7EBF7FBFD7EBF7FBFDFEFF5F9FD7",
            INIT_RAM_37 => X"E773F9DCFEBF3FBFCFE36DB5DAED769B4D9ECF67AFB85C6E171D85AAD12492489C922944",
            INIT_RAM_38 => X"EBF5FAFD7EBF5F9FD7E7F3FAFCFE7F3F9FC7E3F1F9FCFE3F1F8FC7E3F1B8FC6E773B8FCF",
            INIT_RAM_39 => X"EBF7FBFDFEFF5FAFD7EBF5FBFD7EFF5FAFDFEBF5FAFDFEFF7FBFDFEFF5FAFDFEBF7FBFDF",
            INIT_RAM_3A => X"B6D12491389C4E594CC2E9B6DE7F3F9FEFF7FBFDFEFF7FBFDFEFF7EBF5FBFD7EBF5FAFDF",
            INIT_RAM_3B => X"E3F1F8FC6E371B6DC6E773F9DB6E773FAFD7EBF3B6DAED769B5D9ECF67B1B85C763B2D95",
            INIT_RAM_3C => X"EBF7FAFD7EFF5FAFD7EBF3FAFD7EBF3FAFCFE7F3F8FCFEBF1F9FCFE7F3F8FC7E3F1F8FC7",
            INIT_RAM_3D => X"EBF7FAFD7EFF5FAFDFEBF5FAFDFEFF5FAFDFEBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FBFDF",
            INIT_RAM_3E => X"D369B2D85C6E5B2D96BED127924924B26955C76DB8DE7F3FBFEFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_3F => X"E7F3F8FC7E3F1F8FC7E3F1F8FB6DB69B6DCEE7F3F6DB6E773F9FD7E7F3F9FC6DB6BB4DA6"
        )
        port map (
            DO => promx9_inst_15_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_15,
            RESET => reset,
            AD => promx9_inst_15_AD_i
        );

    promx9_inst_16: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"5CAE572B95C9E172B93C1E172783C1E0F0783C1E0F0783C1E0F0373C1E0F0783C1E0F037",
            INIT_RAM_01 => X"DF6FB7DBEDF6FB7DBE7D2E5F4FA5CAE572B95CAE572B93C2E572B95CAE572B93C2E572B8",
            INIT_RAM_02 => X"5CAE4F1F7DA5CE64B158AC0DFECF60B960B1D6695BE1C0E382446817CCFEF3B9EEFB7DBE",
            INIT_RAM_03 => X"3C1E0F0783C0DCF0783C1E0F0373C0DC6E371B8DFEDB558CCB6DF71C0E3EFB5FB8E172FB",
            INIT_RAM_04 => X"5CAE572FA5CAE572FA5CAE1F4B95CAE572B95CAE572B93C2E4F0783C1E172783C1E0F078",
            INIT_RAM_05 => X"17CD4713B9EEFB7DBEDF6FB7DBEDF6FB7DBE5CBE972FA5CBE972FA5CAE572B95CBE9F4B9",
            INIT_RAM_06 => X"3C1E3EFB6FB8E172B97D9E17278FBEDAE8F158BC0DE6FF60BD60B1172A53C1A0F5884A68",
            INIT_RAM_07 => X"3C2E4F0783C1E172783C1E0F0783C1E0F0781C1E0F0783C1E06E781B9E3ED33996D7EE38",
            INIT_RAM_08 => X"7D3E972FA5CAE5F4B95CAE572B97D2E1F4B97D3E972B95CAE572B95CAE572B95CAE572B9",
            INIT_RAM_09 => X"D6DB13DDA4F6904CA917CD5733D9EEFB7DBEDF6FB7DBEDF6FB7DBE5CBE9F4FA5CBE9F4B9",
            INIT_RAM_0A => X"3C0DFED74DB0E0F0783C2E7EFB61B9E1F6B93C7DC70B95CFDF6933783C5606F171BD60B1",
            INIT_RAM_0B => X"5CAE572B95C9E172B93C1E0F0B93C2E4F0785C9E0F0783C1E0F0783C1E0F0383C1E06E78",
            INIT_RAM_0C => X"5CAE5F4B95CBE972B95CBE970FA5CAE572B87D2E572B97D2E5F4B97D2E172FA5CAE572B9",
            INIT_RAM_0D => X"B9BC5E0B0171BD62B137EB5BFDA0F095532AD6ED9F73DBE4F77DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_0E => X"1B9E06E371B8DC6E37FB0DFEDF6FB9E172B93C1E3EFF71C1E0F078FBCD76AB97D9E06D74",
            INIT_RAM_0F => X"5CBE972B95CAE570B95CAE572785C1E0F0785C9E0F0783C1E0F0783C1E0F0783C1E0F078",
            INIT_RAM_10 => X"DF6FB7DBEDF6FB7DBE7D2E172FA5CAE5F4B95CBE972B95CBE972B85CBE970B95CAE1F4B8",
            INIT_RAM_11 => X"99AC66AB97DAE471F7DACCA64B0582C5E2B1580BDC1DA2F19A55ADD6ED5F73B9EEFB7DBE",
            INIT_RAM_12 => X"3C1E0F0783C0DCF0373C0DC6E371BFD86FF61BFD86FF61C0E172783C2E7EFF71B8E071F7",
            INIT_RAM_13 => X"5C9E0F0B95CAE4F0B95CAE170B85C9E0F0785C1E0F0783C2E4F0783C1E0F0783C1E0F078",
            INIT_RAM_14 => X"D6ED6773D9EEFB7DBEDF6FB7DBEDF6FB7DBE5C9E172B93C2E570B95C1E0F0783C1E0F078",
            INIT_RAM_15 => X"1C0DFEFB5FBFDFEF3358CCF6CB97DBED7278FBDD266B1582C162B158AC449DA2F2A2D5AD",
            INIT_RAM_16 => X"3C1E172B93C1E0F0783C1E0F0783C1E0F0783C1E06E781B8DFEC37FB0DC7037FBFDC7038",
            INIT_RAM_17 => X"5CBE972B95CAE5F4B95CAE570B95CAE572B95CAE572785CAE572B93C2E572785CAE57278",
            INIT_RAM_18 => X"58AC551984F3A3582F17FD9F53DBE6FB7DBEDF6FB7DBEDF6FB7DBE7D2E570B95CAE5F4B9",
            INIT_RAM_19 => X"3C0DC7037FBEDB6DB6DB7DF6D74DB6DA66B199EDA6A787DBEDF6B91C6DAE8F1783C56333",
            INIT_RAM_1A => X"5CAE572B95CAE572B85CAE572783C2E572783C1E0F0783C1E0F0783C1E0F0781B9E0F078",
            INIT_RAM_1B => X"5CAE5F4FA5CBE972B97D2E1F4B87D2E570B95CAE5F4B95C3E970B95CAE572B95CAE572B9",
            INIT_RAM_1C => X"5CFDE6AF1782C5633399BC759982E4A45C2E17FDA773DBE6FB7DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_1D => X"3C1E0F0781B9E06E371B8DC7037FBDD3693599CCD6333DA4CE673399FDF6C387DBEDF6FB",
            INIT_RAM_1E => X"5CAE5F4B95CAE572FA5CAE572B95CAE572B95CAE570B93C1E172783C1E0F0783C1E0F078",
            INIT_RAM_1F => X"DF6FB7DBEDF6FB7DBE7D2E572FA5C3E972B97D2E572B97D2E5F4B85CAE572B95CBE972B9",
            INIT_RAM_20 => X"DB7DFEFF75CBEDF6FB5C8DEE93378BC6673399CC85BDA6FDA85A2F380DE777CDF6FB7DBE",
            INIT_RAM_21 => X"3C0E06C381C0E06E371B0DC6C371B0DC6C371B9E07037DB5D266B1583C560B199CCE67B4",
            INIT_RAM_22 => X"5C9E0F0785C1E0F0783C1E170783C1E0F0785C1E0F0B81C0E0F0383C1E0F0783C1E07038",
            INIT_RAM_23 => X"581E2773DBE6FB7DBEDF6FB7DBEDF6FB7DBE5CAE170B93C2E572785C9E0F0785C9E0F078",
            INIT_RAM_24 => X"379BCDE6F99CD76DF6FBFDFEFF73C2E572FB5C8DEE93358BC6653399CCCDE9E2E6B05CB1",
            INIT_RAM_25 => X"1A8D46DF61AFD86BF61AFD86BB41A8D46BB41AFDB6DB6DA6D36A373C0E07037FBCD664B0",
            INIT_RAM_26 => X"3C1E0F0383C1E0F0781B9E0F0381C0E0F0361B0D86C361B0D86C361B0D86C361B0D86DF6",
            INIT_RAM_27 => X"BA4CD61208F7B160B1589E2773DDF6FB7DBEDF6FB7DBEDF6FB7DBE1B1E0F0363C1D8F036",
            INIT_RAM_28 => X"3C0E071B6DB5D266B0378B8DEB1DB6DBEFF71C7DFEDF6FB7DD72FB5C8E36D7458CCA6774",
            INIT_RAM_29 => X"DB6DB6DB6DB6DB6DB6DA6DB69B6DB6DB69B4DA6D2E574DA5CAE9B4B95CAE572B9DCF6A78",
            INIT_RAM_2A => X"1B7D86C351B0D86E371B8DFEDF6FB7DBEDF6FB7DBEDF6FB7DBEDB6FB7DB6DF6DB7DBEDF6",
            INIT_RAM_2B => X"5C8E36D74994CA653399CCDE1E4D22C1633299AE6777C9EEFB7DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_2C => X"995CA6532B94CFEE783C0E06FF7DB4D666F1581B9E1B6FB8E06E371C7DFED35FB7DD72FA",
            INIT_RAM_2D => X"DA6D369B4DA6D2E7B4B9ED369B4B9DCEE7B4DA6D2E773B9DCEE972B95CAE572B95CA6572",
            INIT_RAM_2E => X"DF6FB7DBEDF6FB7DBEDA0D769F6DB6DBEDB4DB6D3EDB61AEDB6DB4DB6DB69B6DA6D369B4",
            INIT_RAM_2F => X"1C7DFEDF71B9E172FA5C8E26B33582C6653399DD1E2A973AC6653399AE67B3DDF6FB7DBE",
            INIT_RAM_30 => X"B95CAE532993C66532784CA64F0995D070783C7DFEFB6DACD666F1582C36DF71B8E07037",
            INIT_RAM_31 => X"FB6D36DB4DA5D36973DA6D369B4DA5CF69B4DA5CEE7B4B9DCEE973B95CEE7B4DA5CAE572",
            INIT_RAM_32 => X"99BEE7B3DDF6FB7DBEDF6FB7DBEDF6FB7DBEDA6D369B6DB0D769B4DB6DB69B4DA6D369B4",
            INIT_RAM_33 => X"78DD06C371C7DC70381C7DF6C383C3ED72B95CFDF6D32582C1E33299CCDE12A174CA6735",
            INIT_RAM_34 => X"BA5CAE772B95CAE572B94CA6572B94CA6532994CA6532996D070381BFDF6DB59ACD66733",
            INIT_RAM_35 => X"DA6D36DB4DA6D36DB4BA6D2E974DA5D2E973B9DCEE7B4DA6D2E7B4B9DCEE973B9DD2E773",
            INIT_RAM_36 => X"58CCD61AC585D2E935BA3EE7B3DDF6FB7DBEDF6FB7DBEDF6FB7DBEDA0D76835DA6DB69F6",
            INIT_RAM_37 => X"1C7DF6DB6BA5CE64B0998E070383C1E0F038FBFD870B95CBEDF4B93C7DF68F0170B8DEB0",
            INIT_RAM_38 => X"B9DCEE772B9DCAE772B95CAE572B94CAE532B94CA657278BC6653278BC664F0BA7DCF078",
            INIT_RAM_39 => X"DA6D369B4DA6D369F6DAEDAE9B4DAED36B74DAED76BB4BA6D369B4BA6D2E974BA5CF69B4",
            INIT_RAM_3A => X"1C0E36870D66B3582E58BCD61AD78DD2E9B4DABEE7B7CDF6FB7DBEDF6FB7DBEDF6FB7DBE",
            INIT_RAM_3B => X"78BC1E372DA0E070381BEDBEFB6DA4CE6732DB0E0F0783C0E07078FB8E0F0FB7DBE9F4FA",
            INIT_RAM_3C => X"BA5D369B4BA6D2E7B4B9DCF6972B9DCAE573B95CE6572B95CAE572994CAE532B94C9E132",
            INIT_RAM_3D => X"DF6FB7DBEDF6FB7DBE1AED36835DA0D769B5DB6DAE9B4DAED36BB5DA6D6E9B5DAED6E974",
            INIT_RAM_3E => X"FBAE572FB7DBE9F4B91C6DA662ED66AB59AC179BCDFAC37DD369B6DB3EA7B3DDF6FB7DBE",
            INIT_RAM_3F => X"995CA6532B93C5E33278CC9E372DB0E0F038FBFDB6DB4DA4CE65B4FB8E0F0783C1E07038"
        )
        port map (
            DO => promx9_inst_16_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_17,
            RESET => reset,
            AD => promx9_inst_16_AD_i
        );

    promx9_inst_17: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"EBF5FAFDFEFF5FBFDFEFF7FAFDFEFF3FAFD7E7F5FAFD7EBF5FAFC7EBF5FAFCFEBF3F9FC7",
            INIT_RAM_01 => X"FBFDFEFF7FBFDFEFF7EBF7FAFD7EFF5FAFDFEBF7FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFDF",
            INIT_RAM_02 => X"EBF5FBFCEE36FB5DA6D369B3D95CAE5B4D96C2D327924924D28955CB6DB9DE7F3FDFEFF7",
            INIT_RAM_03 => X"EBF5FAFD7EBF1FAFD7E7F5F9FC7EBF1F8FC7E3F1F8DB6D36BB8DCEE7F3F9DB6E773FAFDF",
            INIT_RAM_04 => X"EBF7FAFD7EBF5FAFD7EBF7FAFD7EBF7FBFDFEFF7FBFDFEBF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_05 => X"CB6DB9FE7F3FDFEFF7FBFDFEFF7FBFDFEFF7EBF5FBFD7EFF5FBFD7EFF5FBFD7EBF5FAFD7",
            INIT_RAM_06 => X"EFF5F9DC6E773FAFD7EFF7FBFD7E771B6DA6D369B3D9ECAE5B4DA6CB5B6692C925129B55",
            INIT_RAM_07 => X"EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E7F5FAFCFEBF5F8FD7E3F3F8DB6D76DB9DCF",
            INIT_RAM_08 => X"EBF5FBFD7EFF7FAFD7EBF5FAFDFEBF7FAFDFEBF5FBFDFEFF7FBFDFEFF7FBFDFEFF5FAFD7",
            INIT_RAM_09 => X"C2DD669239A512AB6DC76DBBFE7F3FDFEFF7FBFDFEFF7FBFDFEFF7EFF5FCFE7EFF9FAFDF",
            INIT_RAM_0A => X"EBF1F8DB6E373FAFD7EBF5F9DC6E3F5FBFD7E7F3B9FDFEBF3B8DB6D769B4D9ECB67B4DA6",
            INIT_RAM_0B => X"EFF7FBFDFEFF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFCFEBF5FAFD7EBF3FAFCFEBF5F8FD7",
            INIT_RAM_0C => X"EFF5FAFD7EFF5FBFDFEFF5FBFD7EFF5FAFDFEBF5FBFD7EBF7FAFDFEBF7FBFE7EFF7FBFDF",
            INIT_RAM_0D => X"DF69B4DA6CF67B4DA6CF616792392536DB75C2F1BBFE7F7F9FEFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_0E => X"E3F5F8FC7E3F1F8FC7E371F8DC6E777FBFDFEFF3F9DCEE7F7F9FCFE76DB6DDFEFF7F9FB6",
            INIT_RAM_0F => X"EBF5FBFDFEFF7FBFDFEFF7FBFDFEFF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7E7F5F9FD7",
            INIT_RAM_10 => X"FBFDFEFF7FBFDFEFF7EBF7FAFD7EBF5FAFD7EBF5FBFD7EBF5FAFDFEFF5FBFD7EBF7FAFDF",
            INIT_RAM_11 => X"DB69B6DDFEFF5F9FCEDB6BB5DA6D369B4DA6D765A692392596FB85C2EDBBFE7F3FDFEFF7",
            INIT_RAM_12 => X"EBF5FAFCFEBF1F9FC7EBF1F8FC7E3F1B8FC6E3F1B8FC6E7F3FAFDFE7F5F9DCEE3F3F9FCE",
            INIT_RAM_13 => X"EBF5FAFD7EBF5FAFDFEBF7FBFDFEFF5FAFD7EFF5FBFD7EFF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_14 => X"C2EDBCFE7F3FDFEFF7FBFDFEFF7FBFDFEFF7EBF5FAFD7EBF5FBFD7EFF5FAFD7EBF5FAFD7",
            INIT_RAM_15 => X"E7F1F9DB6E773B9DB6D36DB8DD7EFF7FBFD7E76DB6DA6D36BB4DA6D369ACB23925970B85",
            INIT_RAM_16 => X"EBF5FAFD7EBF5FAFD7EBF3FAFD7EBF5F9FD7E7F5F8FD7E3F1F8DC7E371F9FC7E773B9FCF",
            INIT_RAM_17 => X"EBF5FAFD7EBF5FAFD7EBF5FBFD7EFF5FAFDFEFF7FAFD7EFF7FBFDFEFF7FBFDFEBF7FAFD7",
            INIT_RAM_18 => X"D369ADB139A5D70B8ECB71BAFE7F7FDFEFF7FBFDFEFF7FBFDFEFF7EBF5FBFDFEBF5FAFD7",
            INIT_RAM_19 => X"E7F1F9FC7E771B8DC6E373B8DB6E371B6DA6DB71B6DDFEFF7FBFD7E7F1B6DA6D369B4DB6",
            INIT_RAM_1A => X"EFF7FBFDFEFF7FBFDFEFF7FAFD7EBF5FAFD7EBF5FAFD7E7F5FAFD7E7F3FAFD7E3F5FAFCF",
            INIT_RAM_1B => X"EBF5FAFD7EBF5FBFD7EBF7FAFDFEBF5FBFD7EBF5FAFD7EFF5FBFDFEBF7FAFD7EBF7FAFDF",
            INIT_RAM_1C => X"EBF3B6DA6D769B4DB6DB69B0B139A5B72D96CB71BCFE7F7FDFEFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_1D => X"E7F5FAFD7E3F3F8FC7E3F1F9FC7E76DB7DB6DB6DB4DB6E36DB4DB6DB73B8DCFEFF7FBFDF",
            INIT_RAM_1E => X"EBF5FAFDFEBF7FAFD7EFF7FBFDFEFF7FBFD7EFF5FBFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_1F => X"FBFDFEFF7FBFDFEFF7F3F5FBFD7EFF5FBFDFEBF5FAFD7EBF5FAFDFEBF5FAFDFEFF5FBFDF",
            INIT_RAM_20 => X"E373B9DCEEBF7FBFDFEBF1F6DB6D369B6DB6DB6BB1D239E6171D96CB71FCFEFFBFDFEFF7",
            INIT_RAM_21 => X"EBF3F9FCFE7F3F8FC7E7F1F9FC7E7F1F9FC7E3F3F9FC7E36DB6DA6D369B5DA6DB6DB6DC6",
            INIT_RAM_22 => X"EBF5FAFD7EFF5FAFD7EBF5FBFD7EBF5FAFD7EFF5FAFDFE7F3FAFCFEFF5FAFD7EBF5F9FCF",
            INIT_RAM_23 => X"D373FCFE7F7FDFEFF7FBFDFEFF7FBFDFEFF7EFF7FBFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7",
            INIT_RAM_24 => X"CF67B3D9EDB6DB8DC6E773B9DCEEFF5FAFDFEBF1F6DB6D369B5DB6DB69B3D349A6173D96",
            INIT_RAM_25 => X"E7F3F9FC6E7F1B9FC6E7F1B9FC6E7F3F9FBEE7F1B8DC6DF6FB6DC7E7F3F9FC7E76DB5DAE",
            INIT_RAM_26 => X"EBF5FAFCFEBF5FAFD7E3F5FAFCFE7F3FAFCFE7F3F9FCFE7F3F9FCFE7F3F9FCFE7F3F9FC6",
            INIT_RAM_27 => X"DB69B5D44A66574DA6D373FCFE7FBFDFEFF7FBFDFEFF7FBFDFEFF7E7F5FAFCFEBF7FAFCF",
            INIT_RAM_28 => X"E7F3F9FC6E36DB6DA6CF65B3DA6E371B9DCEE7F3B8DC6E373BAFDFEBF3F8DB6D36BB6DB6",
            INIT_RAM_29 => X"E371B8DC6E371B8DC6E371B7DC6E371B7DBEDF6FB6DB6DF6DB6DBEDB6DB6DB6DF6FB6DD7",
            INIT_RAM_2A => X"E7F1B9FCFE7F3F8FC7E3F1F8DC6E371B8DC6E371B8DC6E371B8DC6E371B8DC6E371B8DC6",
            INIT_RAM_2B => X"EFF3F8DB6D76BB5DB6DB6DB4D54AA69B4DAEDB75FCFEFF3FDFEFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_2C => X"D76FB5DAEDB6DB9DDFE7F3F8FCEE36DB6DA6D367B4DC6E773F8FC7E7F3B8DB6E373BBFD7",
            INIT_RAM_2D => X"DF6FB7DBEDF6FB7DBEDF6FB7DBEDF6FB7DBEDF6FB7DBEDF6FB6DB6DB6DB6DB6DB6DB5DB6",
            INIT_RAM_2E => X"FBFDFEFF7FBFDFEFF7E373F8DC6E371B8DBEE371B8DC6E7F1B8DBEE371B8DC6DF6FB7DBE",
            INIT_RAM_2F => X"E7F3B8DCEE3F5FBFD7EBF3F6DB6D769B5DB6DB6DB4D6DBAE9B5DB6DB75FCFE7FBFDFEFF7",
            INIT_RAM_30 => X"DB6DB6DAED769B5DAED76BB5DAED76DB9FD7EBF3B9DC6DB6DB6DA6D369B8DCEE3F3F9FC7",
            INIT_RAM_31 => X"E36FB8DBEDF6DB7DBEDF6FB7DBEDF6FB7DBEDF6FB7DBEDF6FB6DBEDB6FB7DBEDF6DB6DB6",
            INIT_RAM_32 => X"DB77FCFE7FBFDFEFF7FBFDFEFF7FBFDFEFF7E36FB8DC6E373F7DBEE371B7DBEE371B8DBE",
            INIT_RAM_33 => X"D36DB9FC7E7F3B9FCFE7F3B8DCFEFF7FBFDFEFF3B8DAED369B4DAEDB6DB4D75CB6BB6DB6",
            INIT_RAM_34 => X"DB6DB7DB6DB6DB6DB6DB6BB5DB6DB6BB5DAED76BB5DAED76FB9FCFE3F3B8DB6DB6DB6DB6",
            INIT_RAM_35 => X"DF6FB8DBEDF6FB8DBEDB6FB6DB6DF6DB6DBEDF6FB7DBEDF6FB7DBEDF6FB6DBEDF6DB7DBE",
            INIT_RAM_36 => X"D36DB5D85D36DB6DB6DB77FCFE7FBFDFEFF7FBFDFEFF7FBFDFEFF7E373F7DCFDF71B7DC6",
            INIT_RAM_37 => X"E7F3B8DC6DB6FB5DAED373F9FCFEBF7F9FCFE771B9FD7EBF7FAFD7EBF3B8DA6CF65B3DA6",
            INIT_RAM_38 => X"DF6FB7DB6DF6DB7DB6DB6DB7DB6DB6BB6DAEDB6BB5DB6D369B5DAED369B5DA6DB73BAFCF",
            INIT_RAM_39 => X"E371B7DC6E36FB7DC6DB71B6DBEDB6FB6DB6DB6DB6DBEDB6FB7DBEDB6FB6DB6DB6FB7DBE",
            INIT_RAM_3A => X"E7F3F7D96CEE173B96D367B5D85D36DB6DBEDB77FCFEFFBFDFEFF7FBFDFEFF7FBFDFEFF7",
            INIT_RAM_3B => X"D36BB4DB6E373F9FCFE3F1B9DC6DF6DB6DAEE373F9FDFEBF3F9FCFE773FBFDFEFF5FAFD7",
            INIT_RAM_3C => X"DB6DB7DBEDB6FB7DBEDF6FB7DB6DF6DB6DBEDB6FB5DB6DB6DB6DB6D76BB6DAEDB6BB5DAE",
            INIT_RAM_3D => X"FBFDFEFF7FBFDFEFF7E7F1B7DCFDF73F7DB6E371B6DC6DB6FB6DB6DF6DB6DB6DB6DB6DB6",
            INIT_RAM_3E => X"E775FBFDFEFF5FAFD7E7F1B6D96C6E370B85CB67B3D85CF6DB8DC6E375FCFE7FBFDFEFF7",
            INIT_RAM_3F => X"D76DB5DAEDB69B4DAED36BB4DB6E373FAFCFE771B8DBEDF6DB5DC6E773FBFCFE7F7F9FCF"
        )
        port map (
            DO => promx9_inst_17_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_17,
            RESET => reset,
            AD => promx9_inst_17_AD_i
        );

    promx9_inst_18: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 18,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"DF5CF7D73DF5CF6D72DB5CB6D72DB5D36D72DF5CF6D72DF5CB6D72DB5CB5D32DB5CB5D32",
            INIT_RAM_01 => X"DB6D77DB4DB6D77DB4DB6D76D74DB6D76DB5DF6D36D35DB5D36D74DF6D37D73DF6D37DB4",
            INIT_RAM_02 => X"DF6D37DB4E36D39E35DF6D37DB4E36DB6DB5E36DB8DB4DB5D38DB4DB4D78DB4DB5D37DB4",
            INIT_RAM_03 => X"DB6D7BEFBF3CF7CF3DFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
            INIT_RAM_04 => X"E78E38DB6D32C71BACC6EAAFB2ABECA2FB2AC6EB32C2ECB0BAFB2ACAFB36D72E36DB8DB6",
            INIT_RAM_05 => X"E79E3BE78EBAE7BE78EBAE79E78E78E39E38E79E3BEB9EFBEFBEFBF3CEFBEFBEFAE79E38",
            INIT_RAM_06 => X"D74CB4CF1D74CB6D72E36DBBE78E79E39E38E78E39DF7E36DB8DB4E36D36D74E36D39E38",
            INIT_RAM_07 => X"DB5CB6D72D74CB6D72DB5CB6D72DB5CB5D32DB5CB5D32DB5CB5D32D74CB5D32D73C35D32",
            INIT_RAM_08 => X"DF6D36DB5DB6D76D74DB5D37DB4DF5CF7D73DB5CB7DB4DB5CB7DB4DB5CB6D72DB5CB6D72",
            INIT_RAM_09 => X"E36DB6DB5E36DB8DB6DB6D76DB5DB5D36DB5DB5D36DB5DF6D36DB5DB5D36D74DB6D76D74",
            INIT_RAM_0A => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDF6D37DB4DF6D38DB4E36D38DB4E36D36DB5",
            INIT_RAM_0B => X"CAFAB2BECCAFB2EB2ACB0BB6D74E36DB9DF7E37DBBEFBF3CF7EFBEFBEFBEFBEFBEFBEFBE",
            INIT_RAM_0C => X"EFAE7AEFAEFBEFBEFBEFBEFBEFBEFAE7AEB9E77DF8DB6CAFB31BAAC6CA6FB2ABECA2FB2A",
            INIT_RAM_0D => X"E78E39DF7E36DB8DB6E36DB6D35E36DBBE78E78E3AEB9EF9E3AEB9EF9E39E38E78E3AE78",
            INIT_RAM_0E => X"DB5CB4CF1DB5CB4CF1DB5CB4CF1D74CB4CF1D74CB4CF1D74CB6D72E77DF9E38EF9E39E78",
            INIT_RAM_0F => X"DF5CF6D72DB5CB6D72DB5CB6D72DB5CB7D73DB5CB6D72DB5CB6D72DB5CB5D32DB5CB5D32",
            INIT_RAM_10 => X"DB6D76DB5DB5D36D74DB6D76DB5DF6D36D74DB6D76D74DB6D77DB4DF6D37DB4DF5CF6D74",
            INIT_RAM_11 => X"DF6D37DB4E78D77DB4E78D77DB4DF6D38DF6E36DB6DB5DB6D78DB4E36DB6DB5E36DB7DB4",
            INIT_RAM_12 => X"E38DFCF3BF3CEFEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
            INIT_RAM_13 => X"E77DF5D32C6EB30B6AC6CA6FB28BECA2FB28C6EAB2BECC2DAAEB2AD33C37DB4E37DB8DF6",
            INIT_RAM_14 => X"EBAE79E78EFAE7BEB9EBAE79E38E78E3AEB9EFAE7BEFBEFBEFCEFAEFBEFBEB9EB9E39E38",
            INIT_RAM_15 => X"D74CB5D32D33C76D33E77DF9E38E79E39E38E78E38E37E77DF8DF6E36DB8DB6E77DFBE78",
            INIT_RAM_16 => X"DB5CB6D72D74CB6D72DB5CB6D72DB5CB6D72D74CB6D72D74CB6D72D33C76D72D74CB5D32",
            INIT_RAM_17 => X"DF6D36DB5DB6D76D74DB5D37DB4DF5CF7DB4DB5CB7D73DF6D36D72DB5CB6D72DB5CB6D72",
            INIT_RAM_18 => X"E36DB8DB6E36DB6DB5E36DB6DB5E36DB7DB4DB6D76D74DF6D36DB5DB5D36D74DB6D76DB5",
            INIT_RAM_19 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDF6D39E35DF6D37DB4DF6D38DF6DF6D38DB6",
            INIT_RAM_1A => X"C2EB30BACC2DAB1BAADF5CB8DF6E38DF8E37E78E3CF3BF3CF7CF3DFBEFBEFBEFBEFBEFBE",
            INIT_RAM_1B => X"EFAE7CF3BF3CEFBEFBEBBEBAEB9EB9E39E38E36DB4CF1C2EB2FB28BECA2EAE7BECA2FB28",
            INIT_RAM_1C => X"EBAE79DF7E78E39DF7E37DB9DF7E78E3AEB9E78E3BEB9EFAE7BEB9E79E3BE78EF9E3BEFB",
            INIT_RAM_1D => X"D74CB6D72D33C76D72D74CB5D32D33C75D32D74CB5D32DB5CB6D72E38DF9E38EF9E39E78",
            INIT_RAM_1E => X"DB5CB6D72DB5CB6D72DB5CB6D72DF5CF6D72DB5CB6D72DB5CB6D72DB5CB5D32DB5CB5D32",
            INIT_RAM_1F => X"E36DB6DB5DF6D36DB5DB5D37DB4DB6D76DB5DF6D36D74DB6D77DB4DB5D37DB4DF6D37DB4",
            INIT_RAM_20 => X"DF6D37DB4DF6D39E35DF6D39E35DF6D38DB6E36DB8DB6E36DB8DB6DB6D77DB4E36DB6DB5",
            INIT_RAM_21 => X"E78E3CF3BF3CF7EFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBE",
            INIT_RAM_22 => X"DB4D76D72CB0BAEAE7BECA2FB28BECA2FB28C6EAB0B6ABECA33C2EDF5CF8E37E78DB8E37",
            INIT_RAM_23 => X"EBAE7BEB9EFAE7BEB9E79E39E38EFAE7BEFBF3BEBCF3BEFBEFAEFAEFAE7AEB9E78E39DF7",
            INIT_RAM_24 => X"D74CB5D32D74CB6D74E38DF9E38E79E3BE78EB9E39E38E77DF8E37E77DF8E37EBAE7BE78",
            INIT_RAM_25 => X"DB5CB6D72DB5CB6D72DB5CB6D72DB5CB6D72D33C76D72D74CB6D72D74CB6D72D74CB5D32",
            INIT_RAM_26 => X"DB5D36DB5DB6D76DB5DB5D37D73DF6D37DB4DB5CB7DB4DB5CB7DB4DB5CB6D72DB5CB6D72",
            INIT_RAM_27 => X"E36DB8DB6DB6D78DB6DB6D78DB6E36DB6DB5E36DB6D74DB5D36DB5DB6D77DB4DB6D76DB5",
            INIT_RAM_28 => X"FBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEFBEDF6D39E35DF6D37DB4DF6D37DB4E36DB6DB5",
            INIT_RAM_29 => X"C2DAB1B29BECAB5D32E36DB8DF6E38DF9E38E78E3CF3BF3CF7EFBEFBEFBEFBEFBEFBEFBE",
            INIT_RAM_2A => X"F3BEBCF3BEFBEFAEFAEFAE7BE78EF9E39DF7DB4CF5D32CF0BAEAE7BAB9EEAE7BECA2FB28",
            INIT_RAM_2B => X"EF9E39E38E77DF9DF7E38DF9E38EF9E3BE78EBAE7BEB9EFAE7BEB9E78E3BEB9EFBEFCEFA",
            INIT_RAM_2C => X"D74CB6D72D74CB5D32D74CB4CF1D74CB5D32D74CB5CF0DB5CB6D72E77DF9E38EF9E39E78",
            INIT_RAM_2D => X"DB5CB6D72DB5CB6D72DB5CB6D72DF5CF6D72DB5CB6D72DB5CB6D72DB5CB5D32DB5CB5D32",
            INIT_RAM_2E => X"E36DB6DB5DB5D36DB5DF6D36D74DB5D36D74DB5D36D74DB5D36D74DB5D37D73DB5CB6D74",
            INIT_RAM_2F => X"DF6D37DB4DF6D39E35E36D39E35DF6D38DB6E36DB8DB6DB6D78DB6DF6D36DB5DB6D77DB4"
        )
        port map (
            DO => promx9_inst_18_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_19,
            RESET => reset,
            AD => promx9_inst_18_AD_i
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ad(14),
            CLK => clk,
            CE => ce
        );

    dff_inst_1: DFFE
        port map (
            Q => dff_q_1,
            D => ad(13),
            CLK => clk,
            CE => ce
        );

    dff_inst_2: DFFE
        port map (
            Q => dff_q_2,
            D => ad(12),
            CLK => clk,
            CE => ce
        );

    dff_inst_3: DFFE
        port map (
            Q => dff_q_3,
            D => ad(11),
            CLK => clk,
            CE => ce
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => promx9_inst_0_dout(0),
            I1 => promx9_inst_1_dout(0),
            S0 => dff_q_3
        );

    mux_inst_11: MUX2
        port map (
            O => mux_o_11,
            I0 => promx9_inst_2_dout(0),
            I1 => promx9_inst_3_dout(0),
            S0 => dff_q_3
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => promx9_inst_4_dout(0),
            I1 => promx9_inst_5_dout(0),
            S0 => dff_q_3
        );

    mux_inst_13: MUX2
        port map (
            O => mux_o_13,
            I0 => promx9_inst_6_dout(0),
            I1 => promx9_inst_7_dout(0),
            S0 => dff_q_3
        );

    mux_inst_14: MUX2
        port map (
            O => mux_o_14,
            I0 => promx9_inst_16_dout(0),
            I1 => promx9_inst_18_dout(0),
            S0 => dff_q_3
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => mux_o_10,
            I1 => mux_o_11,
            S0 => dff_q_2
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => mux_o_12,
            I1 => mux_o_13,
            S0 => dff_q_2
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => mux_o_15,
            I1 => mux_o_16,
            S0 => dff_q_1
        );

    mux_inst_20: MUX2
        port map (
            O => dout(0),
            I0 => mux_o_18,
            I1 => mux_o_14,
            S0 => dff_q_0
        );

    mux_inst_31: MUX2
        port map (
            O => mux_o_31,
            I0 => promx9_inst_0_dout(1),
            I1 => promx9_inst_1_dout(1),
            S0 => dff_q_3
        );

    mux_inst_32: MUX2
        port map (
            O => mux_o_32,
            I0 => promx9_inst_2_dout(1),
            I1 => promx9_inst_3_dout(1),
            S0 => dff_q_3
        );

    mux_inst_33: MUX2
        port map (
            O => mux_o_33,
            I0 => promx9_inst_4_dout(1),
            I1 => promx9_inst_5_dout(1),
            S0 => dff_q_3
        );

    mux_inst_34: MUX2
        port map (
            O => mux_o_34,
            I0 => promx9_inst_6_dout(1),
            I1 => promx9_inst_7_dout(1),
            S0 => dff_q_3
        );

    mux_inst_35: MUX2
        port map (
            O => mux_o_35,
            I0 => promx9_inst_16_dout(1),
            I1 => promx9_inst_18_dout(1),
            S0 => dff_q_3
        );

    mux_inst_36: MUX2
        port map (
            O => mux_o_36,
            I0 => mux_o_31,
            I1 => mux_o_32,
            S0 => dff_q_2
        );

    mux_inst_37: MUX2
        port map (
            O => mux_o_37,
            I0 => mux_o_33,
            I1 => mux_o_34,
            S0 => dff_q_2
        );

    mux_inst_39: MUX2
        port map (
            O => mux_o_39,
            I0 => mux_o_36,
            I1 => mux_o_37,
            S0 => dff_q_1
        );

    mux_inst_41: MUX2
        port map (
            O => dout(1),
            I0 => mux_o_39,
            I1 => mux_o_35,
            S0 => dff_q_0
        );

    mux_inst_52: MUX2
        port map (
            O => mux_o_52,
            I0 => promx9_inst_0_dout(2),
            I1 => promx9_inst_1_dout(2),
            S0 => dff_q_3
        );

    mux_inst_53: MUX2
        port map (
            O => mux_o_53,
            I0 => promx9_inst_2_dout(2),
            I1 => promx9_inst_3_dout(2),
            S0 => dff_q_3
        );

    mux_inst_54: MUX2
        port map (
            O => mux_o_54,
            I0 => promx9_inst_4_dout(2),
            I1 => promx9_inst_5_dout(2),
            S0 => dff_q_3
        );

    mux_inst_55: MUX2
        port map (
            O => mux_o_55,
            I0 => promx9_inst_6_dout(2),
            I1 => promx9_inst_7_dout(2),
            S0 => dff_q_3
        );

    mux_inst_56: MUX2
        port map (
            O => mux_o_56,
            I0 => promx9_inst_16_dout(2),
            I1 => promx9_inst_18_dout(2),
            S0 => dff_q_3
        );

    mux_inst_57: MUX2
        port map (
            O => mux_o_57,
            I0 => mux_o_52,
            I1 => mux_o_53,
            S0 => dff_q_2
        );

    mux_inst_58: MUX2
        port map (
            O => mux_o_58,
            I0 => mux_o_54,
            I1 => mux_o_55,
            S0 => dff_q_2
        );

    mux_inst_60: MUX2
        port map (
            O => mux_o_60,
            I0 => mux_o_57,
            I1 => mux_o_58,
            S0 => dff_q_1
        );

    mux_inst_62: MUX2
        port map (
            O => dout(2),
            I0 => mux_o_60,
            I1 => mux_o_56,
            S0 => dff_q_0
        );

    mux_inst_73: MUX2
        port map (
            O => mux_o_73,
            I0 => promx9_inst_0_dout(3),
            I1 => promx9_inst_1_dout(3),
            S0 => dff_q_3
        );

    mux_inst_74: MUX2
        port map (
            O => mux_o_74,
            I0 => promx9_inst_2_dout(3),
            I1 => promx9_inst_3_dout(3),
            S0 => dff_q_3
        );

    mux_inst_75: MUX2
        port map (
            O => mux_o_75,
            I0 => promx9_inst_4_dout(3),
            I1 => promx9_inst_5_dout(3),
            S0 => dff_q_3
        );

    mux_inst_76: MUX2
        port map (
            O => mux_o_76,
            I0 => promx9_inst_6_dout(3),
            I1 => promx9_inst_7_dout(3),
            S0 => dff_q_3
        );

    mux_inst_77: MUX2
        port map (
            O => mux_o_77,
            I0 => promx9_inst_16_dout(3),
            I1 => promx9_inst_18_dout(3),
            S0 => dff_q_3
        );

    mux_inst_78: MUX2
        port map (
            O => mux_o_78,
            I0 => mux_o_73,
            I1 => mux_o_74,
            S0 => dff_q_2
        );

    mux_inst_79: MUX2
        port map (
            O => mux_o_79,
            I0 => mux_o_75,
            I1 => mux_o_76,
            S0 => dff_q_2
        );

    mux_inst_81: MUX2
        port map (
            O => mux_o_81,
            I0 => mux_o_78,
            I1 => mux_o_79,
            S0 => dff_q_1
        );

    mux_inst_83: MUX2
        port map (
            O => dout(3),
            I0 => mux_o_81,
            I1 => mux_o_77,
            S0 => dff_q_0
        );

    mux_inst_94: MUX2
        port map (
            O => mux_o_94,
            I0 => promx9_inst_0_dout(4),
            I1 => promx9_inst_1_dout(4),
            S0 => dff_q_3
        );

    mux_inst_95: MUX2
        port map (
            O => mux_o_95,
            I0 => promx9_inst_2_dout(4),
            I1 => promx9_inst_3_dout(4),
            S0 => dff_q_3
        );

    mux_inst_96: MUX2
        port map (
            O => mux_o_96,
            I0 => promx9_inst_4_dout(4),
            I1 => promx9_inst_5_dout(4),
            S0 => dff_q_3
        );

    mux_inst_97: MUX2
        port map (
            O => mux_o_97,
            I0 => promx9_inst_6_dout(4),
            I1 => promx9_inst_7_dout(4),
            S0 => dff_q_3
        );

    mux_inst_98: MUX2
        port map (
            O => mux_o_98,
            I0 => promx9_inst_16_dout(4),
            I1 => promx9_inst_18_dout(4),
            S0 => dff_q_3
        );

    mux_inst_99: MUX2
        port map (
            O => mux_o_99,
            I0 => mux_o_94,
            I1 => mux_o_95,
            S0 => dff_q_2
        );

    mux_inst_100: MUX2
        port map (
            O => mux_o_100,
            I0 => mux_o_96,
            I1 => mux_o_97,
            S0 => dff_q_2
        );

    mux_inst_102: MUX2
        port map (
            O => mux_o_102,
            I0 => mux_o_99,
            I1 => mux_o_100,
            S0 => dff_q_1
        );

    mux_inst_104: MUX2
        port map (
            O => dout(4),
            I0 => mux_o_102,
            I1 => mux_o_98,
            S0 => dff_q_0
        );

    mux_inst_115: MUX2
        port map (
            O => mux_o_115,
            I0 => promx9_inst_0_dout(5),
            I1 => promx9_inst_1_dout(5),
            S0 => dff_q_3
        );

    mux_inst_116: MUX2
        port map (
            O => mux_o_116,
            I0 => promx9_inst_2_dout(5),
            I1 => promx9_inst_3_dout(5),
            S0 => dff_q_3
        );

    mux_inst_117: MUX2
        port map (
            O => mux_o_117,
            I0 => promx9_inst_4_dout(5),
            I1 => promx9_inst_5_dout(5),
            S0 => dff_q_3
        );

    mux_inst_118: MUX2
        port map (
            O => mux_o_118,
            I0 => promx9_inst_6_dout(5),
            I1 => promx9_inst_7_dout(5),
            S0 => dff_q_3
        );

    mux_inst_119: MUX2
        port map (
            O => mux_o_119,
            I0 => promx9_inst_16_dout(5),
            I1 => promx9_inst_18_dout(5),
            S0 => dff_q_3
        );

    mux_inst_120: MUX2
        port map (
            O => mux_o_120,
            I0 => mux_o_115,
            I1 => mux_o_116,
            S0 => dff_q_2
        );

    mux_inst_121: MUX2
        port map (
            O => mux_o_121,
            I0 => mux_o_117,
            I1 => mux_o_118,
            S0 => dff_q_2
        );

    mux_inst_123: MUX2
        port map (
            O => mux_o_123,
            I0 => mux_o_120,
            I1 => mux_o_121,
            S0 => dff_q_1
        );

    mux_inst_125: MUX2
        port map (
            O => dout(5),
            I0 => mux_o_123,
            I1 => mux_o_119,
            S0 => dff_q_0
        );

    mux_inst_136: MUX2
        port map (
            O => mux_o_136,
            I0 => promx9_inst_0_dout(6),
            I1 => promx9_inst_1_dout(6),
            S0 => dff_q_3
        );

    mux_inst_137: MUX2
        port map (
            O => mux_o_137,
            I0 => promx9_inst_2_dout(6),
            I1 => promx9_inst_3_dout(6),
            S0 => dff_q_3
        );

    mux_inst_138: MUX2
        port map (
            O => mux_o_138,
            I0 => promx9_inst_4_dout(6),
            I1 => promx9_inst_5_dout(6),
            S0 => dff_q_3
        );

    mux_inst_139: MUX2
        port map (
            O => mux_o_139,
            I0 => promx9_inst_6_dout(6),
            I1 => promx9_inst_7_dout(6),
            S0 => dff_q_3
        );

    mux_inst_140: MUX2
        port map (
            O => mux_o_140,
            I0 => promx9_inst_16_dout(6),
            I1 => promx9_inst_18_dout(6),
            S0 => dff_q_3
        );

    mux_inst_141: MUX2
        port map (
            O => mux_o_141,
            I0 => mux_o_136,
            I1 => mux_o_137,
            S0 => dff_q_2
        );

    mux_inst_142: MUX2
        port map (
            O => mux_o_142,
            I0 => mux_o_138,
            I1 => mux_o_139,
            S0 => dff_q_2
        );

    mux_inst_144: MUX2
        port map (
            O => mux_o_144,
            I0 => mux_o_141,
            I1 => mux_o_142,
            S0 => dff_q_1
        );

    mux_inst_146: MUX2
        port map (
            O => dout(6),
            I0 => mux_o_144,
            I1 => mux_o_140,
            S0 => dff_q_0
        );

    mux_inst_157: MUX2
        port map (
            O => mux_o_157,
            I0 => promx9_inst_0_dout(7),
            I1 => promx9_inst_1_dout(7),
            S0 => dff_q_3
        );

    mux_inst_158: MUX2
        port map (
            O => mux_o_158,
            I0 => promx9_inst_2_dout(7),
            I1 => promx9_inst_3_dout(7),
            S0 => dff_q_3
        );

    mux_inst_159: MUX2
        port map (
            O => mux_o_159,
            I0 => promx9_inst_4_dout(7),
            I1 => promx9_inst_5_dout(7),
            S0 => dff_q_3
        );

    mux_inst_160: MUX2
        port map (
            O => mux_o_160,
            I0 => promx9_inst_6_dout(7),
            I1 => promx9_inst_7_dout(7),
            S0 => dff_q_3
        );

    mux_inst_161: MUX2
        port map (
            O => mux_o_161,
            I0 => promx9_inst_16_dout(7),
            I1 => promx9_inst_18_dout(7),
            S0 => dff_q_3
        );

    mux_inst_162: MUX2
        port map (
            O => mux_o_162,
            I0 => mux_o_157,
            I1 => mux_o_158,
            S0 => dff_q_2
        );

    mux_inst_163: MUX2
        port map (
            O => mux_o_163,
            I0 => mux_o_159,
            I1 => mux_o_160,
            S0 => dff_q_2
        );

    mux_inst_165: MUX2
        port map (
            O => mux_o_165,
            I0 => mux_o_162,
            I1 => mux_o_163,
            S0 => dff_q_1
        );

    mux_inst_167: MUX2
        port map (
            O => dout(7),
            I0 => mux_o_165,
            I1 => mux_o_161,
            S0 => dff_q_0
        );

    mux_inst_178: MUX2
        port map (
            O => mux_o_178,
            I0 => promx9_inst_0_dout(8),
            I1 => promx9_inst_1_dout(8),
            S0 => dff_q_3
        );

    mux_inst_179: MUX2
        port map (
            O => mux_o_179,
            I0 => promx9_inst_2_dout(8),
            I1 => promx9_inst_3_dout(8),
            S0 => dff_q_3
        );

    mux_inst_180: MUX2
        port map (
            O => mux_o_180,
            I0 => promx9_inst_4_dout(8),
            I1 => promx9_inst_5_dout(8),
            S0 => dff_q_3
        );

    mux_inst_181: MUX2
        port map (
            O => mux_o_181,
            I0 => promx9_inst_6_dout(8),
            I1 => promx9_inst_7_dout(8),
            S0 => dff_q_3
        );

    mux_inst_182: MUX2
        port map (
            O => mux_o_182,
            I0 => promx9_inst_16_dout(8),
            I1 => promx9_inst_18_dout(8),
            S0 => dff_q_3
        );

    mux_inst_183: MUX2
        port map (
            O => mux_o_183,
            I0 => mux_o_178,
            I1 => mux_o_179,
            S0 => dff_q_2
        );

    mux_inst_184: MUX2
        port map (
            O => mux_o_184,
            I0 => mux_o_180,
            I1 => mux_o_181,
            S0 => dff_q_2
        );

    mux_inst_186: MUX2
        port map (
            O => mux_o_186,
            I0 => mux_o_183,
            I1 => mux_o_184,
            S0 => dff_q_1
        );

    mux_inst_188: MUX2
        port map (
            O => dout(8),
            I0 => mux_o_186,
            I1 => mux_o_182,
            S0 => dff_q_0
        );

    mux_inst_199: MUX2
        port map (
            O => mux_o_199,
            I0 => promx9_inst_8_dout(9),
            I1 => promx9_inst_9_dout(9),
            S0 => dff_q_3
        );

    mux_inst_200: MUX2
        port map (
            O => mux_o_200,
            I0 => promx9_inst_10_dout(9),
            I1 => promx9_inst_11_dout(9),
            S0 => dff_q_3
        );

    mux_inst_201: MUX2
        port map (
            O => mux_o_201,
            I0 => promx9_inst_12_dout(9),
            I1 => promx9_inst_13_dout(9),
            S0 => dff_q_3
        );

    mux_inst_202: MUX2
        port map (
            O => mux_o_202,
            I0 => promx9_inst_14_dout(9),
            I1 => promx9_inst_15_dout(9),
            S0 => dff_q_3
        );

    mux_inst_203: MUX2
        port map (
            O => mux_o_203,
            I0 => promx9_inst_17_dout(9),
            I1 => promx9_inst_18_dout(9),
            S0 => dff_q_3
        );

    mux_inst_204: MUX2
        port map (
            O => mux_o_204,
            I0 => mux_o_199,
            I1 => mux_o_200,
            S0 => dff_q_2
        );

    mux_inst_205: MUX2
        port map (
            O => mux_o_205,
            I0 => mux_o_201,
            I1 => mux_o_202,
            S0 => dff_q_2
        );

    mux_inst_207: MUX2
        port map (
            O => mux_o_207,
            I0 => mux_o_204,
            I1 => mux_o_205,
            S0 => dff_q_1
        );

    mux_inst_209: MUX2
        port map (
            O => dout(9),
            I0 => mux_o_207,
            I1 => mux_o_203,
            S0 => dff_q_0
        );

    mux_inst_220: MUX2
        port map (
            O => mux_o_220,
            I0 => promx9_inst_8_dout(10),
            I1 => promx9_inst_9_dout(10),
            S0 => dff_q_3
        );

    mux_inst_221: MUX2
        port map (
            O => mux_o_221,
            I0 => promx9_inst_10_dout(10),
            I1 => promx9_inst_11_dout(10),
            S0 => dff_q_3
        );

    mux_inst_222: MUX2
        port map (
            O => mux_o_222,
            I0 => promx9_inst_12_dout(10),
            I1 => promx9_inst_13_dout(10),
            S0 => dff_q_3
        );

    mux_inst_223: MUX2
        port map (
            O => mux_o_223,
            I0 => promx9_inst_14_dout(10),
            I1 => promx9_inst_15_dout(10),
            S0 => dff_q_3
        );

    mux_inst_224: MUX2
        port map (
            O => mux_o_224,
            I0 => promx9_inst_17_dout(10),
            I1 => promx9_inst_18_dout(10),
            S0 => dff_q_3
        );

    mux_inst_225: MUX2
        port map (
            O => mux_o_225,
            I0 => mux_o_220,
            I1 => mux_o_221,
            S0 => dff_q_2
        );

    mux_inst_226: MUX2
        port map (
            O => mux_o_226,
            I0 => mux_o_222,
            I1 => mux_o_223,
            S0 => dff_q_2
        );

    mux_inst_228: MUX2
        port map (
            O => mux_o_228,
            I0 => mux_o_225,
            I1 => mux_o_226,
            S0 => dff_q_1
        );

    mux_inst_230: MUX2
        port map (
            O => dout(10),
            I0 => mux_o_228,
            I1 => mux_o_224,
            S0 => dff_q_0
        );

    mux_inst_241: MUX2
        port map (
            O => mux_o_241,
            I0 => promx9_inst_8_dout(11),
            I1 => promx9_inst_9_dout(11),
            S0 => dff_q_3
        );

    mux_inst_242: MUX2
        port map (
            O => mux_o_242,
            I0 => promx9_inst_10_dout(11),
            I1 => promx9_inst_11_dout(11),
            S0 => dff_q_3
        );

    mux_inst_243: MUX2
        port map (
            O => mux_o_243,
            I0 => promx9_inst_12_dout(11),
            I1 => promx9_inst_13_dout(11),
            S0 => dff_q_3
        );

    mux_inst_244: MUX2
        port map (
            O => mux_o_244,
            I0 => promx9_inst_14_dout(11),
            I1 => promx9_inst_15_dout(11),
            S0 => dff_q_3
        );

    mux_inst_245: MUX2
        port map (
            O => mux_o_245,
            I0 => promx9_inst_17_dout(11),
            I1 => promx9_inst_18_dout(11),
            S0 => dff_q_3
        );

    mux_inst_246: MUX2
        port map (
            O => mux_o_246,
            I0 => mux_o_241,
            I1 => mux_o_242,
            S0 => dff_q_2
        );

    mux_inst_247: MUX2
        port map (
            O => mux_o_247,
            I0 => mux_o_243,
            I1 => mux_o_244,
            S0 => dff_q_2
        );

    mux_inst_249: MUX2
        port map (
            O => mux_o_249,
            I0 => mux_o_246,
            I1 => mux_o_247,
            S0 => dff_q_1
        );

    mux_inst_251: MUX2
        port map (
            O => dout(11),
            I0 => mux_o_249,
            I1 => mux_o_245,
            S0 => dff_q_0
        );

    mux_inst_262: MUX2
        port map (
            O => mux_o_262,
            I0 => promx9_inst_8_dout(12),
            I1 => promx9_inst_9_dout(12),
            S0 => dff_q_3
        );

    mux_inst_263: MUX2
        port map (
            O => mux_o_263,
            I0 => promx9_inst_10_dout(12),
            I1 => promx9_inst_11_dout(12),
            S0 => dff_q_3
        );

    mux_inst_264: MUX2
        port map (
            O => mux_o_264,
            I0 => promx9_inst_12_dout(12),
            I1 => promx9_inst_13_dout(12),
            S0 => dff_q_3
        );

    mux_inst_265: MUX2
        port map (
            O => mux_o_265,
            I0 => promx9_inst_14_dout(12),
            I1 => promx9_inst_15_dout(12),
            S0 => dff_q_3
        );

    mux_inst_266: MUX2
        port map (
            O => mux_o_266,
            I0 => promx9_inst_17_dout(12),
            I1 => promx9_inst_18_dout(12),
            S0 => dff_q_3
        );

    mux_inst_267: MUX2
        port map (
            O => mux_o_267,
            I0 => mux_o_262,
            I1 => mux_o_263,
            S0 => dff_q_2
        );

    mux_inst_268: MUX2
        port map (
            O => mux_o_268,
            I0 => mux_o_264,
            I1 => mux_o_265,
            S0 => dff_q_2
        );

    mux_inst_270: MUX2
        port map (
            O => mux_o_270,
            I0 => mux_o_267,
            I1 => mux_o_268,
            S0 => dff_q_1
        );

    mux_inst_272: MUX2
        port map (
            O => dout(12),
            I0 => mux_o_270,
            I1 => mux_o_266,
            S0 => dff_q_0
        );

    mux_inst_283: MUX2
        port map (
            O => mux_o_283,
            I0 => promx9_inst_8_dout(13),
            I1 => promx9_inst_9_dout(13),
            S0 => dff_q_3
        );

    mux_inst_284: MUX2
        port map (
            O => mux_o_284,
            I0 => promx9_inst_10_dout(13),
            I1 => promx9_inst_11_dout(13),
            S0 => dff_q_3
        );

    mux_inst_285: MUX2
        port map (
            O => mux_o_285,
            I0 => promx9_inst_12_dout(13),
            I1 => promx9_inst_13_dout(13),
            S0 => dff_q_3
        );

    mux_inst_286: MUX2
        port map (
            O => mux_o_286,
            I0 => promx9_inst_14_dout(13),
            I1 => promx9_inst_15_dout(13),
            S0 => dff_q_3
        );

    mux_inst_287: MUX2
        port map (
            O => mux_o_287,
            I0 => promx9_inst_17_dout(13),
            I1 => promx9_inst_18_dout(13),
            S0 => dff_q_3
        );

    mux_inst_288: MUX2
        port map (
            O => mux_o_288,
            I0 => mux_o_283,
            I1 => mux_o_284,
            S0 => dff_q_2
        );

    mux_inst_289: MUX2
        port map (
            O => mux_o_289,
            I0 => mux_o_285,
            I1 => mux_o_286,
            S0 => dff_q_2
        );

    mux_inst_291: MUX2
        port map (
            O => mux_o_291,
            I0 => mux_o_288,
            I1 => mux_o_289,
            S0 => dff_q_1
        );

    mux_inst_293: MUX2
        port map (
            O => dout(13),
            I0 => mux_o_291,
            I1 => mux_o_287,
            S0 => dff_q_0
        );

    mux_inst_304: MUX2
        port map (
            O => mux_o_304,
            I0 => promx9_inst_8_dout(14),
            I1 => promx9_inst_9_dout(14),
            S0 => dff_q_3
        );

    mux_inst_305: MUX2
        port map (
            O => mux_o_305,
            I0 => promx9_inst_10_dout(14),
            I1 => promx9_inst_11_dout(14),
            S0 => dff_q_3
        );

    mux_inst_306: MUX2
        port map (
            O => mux_o_306,
            I0 => promx9_inst_12_dout(14),
            I1 => promx9_inst_13_dout(14),
            S0 => dff_q_3
        );

    mux_inst_307: MUX2
        port map (
            O => mux_o_307,
            I0 => promx9_inst_14_dout(14),
            I1 => promx9_inst_15_dout(14),
            S0 => dff_q_3
        );

    mux_inst_308: MUX2
        port map (
            O => mux_o_308,
            I0 => promx9_inst_17_dout(14),
            I1 => promx9_inst_18_dout(14),
            S0 => dff_q_3
        );

    mux_inst_309: MUX2
        port map (
            O => mux_o_309,
            I0 => mux_o_304,
            I1 => mux_o_305,
            S0 => dff_q_2
        );

    mux_inst_310: MUX2
        port map (
            O => mux_o_310,
            I0 => mux_o_306,
            I1 => mux_o_307,
            S0 => dff_q_2
        );

    mux_inst_312: MUX2
        port map (
            O => mux_o_312,
            I0 => mux_o_309,
            I1 => mux_o_310,
            S0 => dff_q_1
        );

    mux_inst_314: MUX2
        port map (
            O => dout(14),
            I0 => mux_o_312,
            I1 => mux_o_308,
            S0 => dff_q_0
        );

    mux_inst_325: MUX2
        port map (
            O => mux_o_325,
            I0 => promx9_inst_8_dout(15),
            I1 => promx9_inst_9_dout(15),
            S0 => dff_q_3
        );

    mux_inst_326: MUX2
        port map (
            O => mux_o_326,
            I0 => promx9_inst_10_dout(15),
            I1 => promx9_inst_11_dout(15),
            S0 => dff_q_3
        );

    mux_inst_327: MUX2
        port map (
            O => mux_o_327,
            I0 => promx9_inst_12_dout(15),
            I1 => promx9_inst_13_dout(15),
            S0 => dff_q_3
        );

    mux_inst_328: MUX2
        port map (
            O => mux_o_328,
            I0 => promx9_inst_14_dout(15),
            I1 => promx9_inst_15_dout(15),
            S0 => dff_q_3
        );

    mux_inst_329: MUX2
        port map (
            O => mux_o_329,
            I0 => promx9_inst_17_dout(15),
            I1 => promx9_inst_18_dout(15),
            S0 => dff_q_3
        );

    mux_inst_330: MUX2
        port map (
            O => mux_o_330,
            I0 => mux_o_325,
            I1 => mux_o_326,
            S0 => dff_q_2
        );

    mux_inst_331: MUX2
        port map (
            O => mux_o_331,
            I0 => mux_o_327,
            I1 => mux_o_328,
            S0 => dff_q_2
        );

    mux_inst_333: MUX2
        port map (
            O => mux_o_333,
            I0 => mux_o_330,
            I1 => mux_o_331,
            S0 => dff_q_1
        );

    mux_inst_335: MUX2
        port map (
            O => dout(15),
            I0 => mux_o_333,
            I1 => mux_o_329,
            S0 => dff_q_0
        );

    mux_inst_346: MUX2
        port map (
            O => mux_o_346,
            I0 => promx9_inst_8_dout(16),
            I1 => promx9_inst_9_dout(16),
            S0 => dff_q_3
        );

    mux_inst_347: MUX2
        port map (
            O => mux_o_347,
            I0 => promx9_inst_10_dout(16),
            I1 => promx9_inst_11_dout(16),
            S0 => dff_q_3
        );

    mux_inst_348: MUX2
        port map (
            O => mux_o_348,
            I0 => promx9_inst_12_dout(16),
            I1 => promx9_inst_13_dout(16),
            S0 => dff_q_3
        );

    mux_inst_349: MUX2
        port map (
            O => mux_o_349,
            I0 => promx9_inst_14_dout(16),
            I1 => promx9_inst_15_dout(16),
            S0 => dff_q_3
        );

    mux_inst_350: MUX2
        port map (
            O => mux_o_350,
            I0 => promx9_inst_17_dout(16),
            I1 => promx9_inst_18_dout(16),
            S0 => dff_q_3
        );

    mux_inst_351: MUX2
        port map (
            O => mux_o_351,
            I0 => mux_o_346,
            I1 => mux_o_347,
            S0 => dff_q_2
        );

    mux_inst_352: MUX2
        port map (
            O => mux_o_352,
            I0 => mux_o_348,
            I1 => mux_o_349,
            S0 => dff_q_2
        );

    mux_inst_354: MUX2
        port map (
            O => mux_o_354,
            I0 => mux_o_351,
            I1 => mux_o_352,
            S0 => dff_q_1
        );

    mux_inst_356: MUX2
        port map (
            O => dout(16),
            I0 => mux_o_354,
            I1 => mux_o_350,
            S0 => dff_q_0
        );

    mux_inst_367: MUX2
        port map (
            O => mux_o_367,
            I0 => promx9_inst_8_dout(17),
            I1 => promx9_inst_9_dout(17),
            S0 => dff_q_3
        );

    mux_inst_368: MUX2
        port map (
            O => mux_o_368,
            I0 => promx9_inst_10_dout(17),
            I1 => promx9_inst_11_dout(17),
            S0 => dff_q_3
        );

    mux_inst_369: MUX2
        port map (
            O => mux_o_369,
            I0 => promx9_inst_12_dout(17),
            I1 => promx9_inst_13_dout(17),
            S0 => dff_q_3
        );

    mux_inst_370: MUX2
        port map (
            O => mux_o_370,
            I0 => promx9_inst_14_dout(17),
            I1 => promx9_inst_15_dout(17),
            S0 => dff_q_3
        );

    mux_inst_371: MUX2
        port map (
            O => mux_o_371,
            I0 => promx9_inst_17_dout(17),
            I1 => promx9_inst_18_dout(17),
            S0 => dff_q_3
        );

    mux_inst_372: MUX2
        port map (
            O => mux_o_372,
            I0 => mux_o_367,
            I1 => mux_o_368,
            S0 => dff_q_2
        );

    mux_inst_373: MUX2
        port map (
            O => mux_o_373,
            I0 => mux_o_369,
            I1 => mux_o_370,
            S0 => dff_q_2
        );

    mux_inst_375: MUX2
        port map (
            O => mux_o_375,
            I0 => mux_o_372,
            I1 => mux_o_373,
            S0 => dff_q_1
        );

    mux_inst_377: MUX2
        port map (
            O => dout(17),
            I0 => mux_o_375,
            I1 => mux_o_371,
            S0 => dff_q_0
        );

end Behavioral; --Gowin_pROM
