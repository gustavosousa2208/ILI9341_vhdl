--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.07
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Thu Dec 15 22:40:54 2022

library IEEE;
use IEEE.std_logic_1164.all;

entity gato_colorido is
    port (
        dout: out std_logic_vector(17 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(14 downto 0)
    );
end gato_colorido;

architecture Behavioral of gato_colorido is

    signal lut_f_0: std_logic;
    signal lut_f_1: std_logic;
    signal lut_f_2: std_logic;
    signal lut_f_3: std_logic;
    signal lut_f_4: std_logic;
    signal lut_f_5: std_logic;
    signal lut_f_6: std_logic;
    signal lut_f_7: std_logic;
    signal lut_f_8: std_logic;
    signal lut_f_9: std_logic;
    signal lut_f_10: std_logic;
    signal lut_f_11: std_logic;
    signal lut_f_12: std_logic;
    signal lut_f_13: std_logic;
    signal lut_f_14: std_logic;
    signal lut_f_15: std_logic;
    signal lut_f_16: std_logic;
    signal lut_f_17: std_logic;
    signal lut_f_18: std_logic;
    signal lut_f_19: std_logic;
    signal promx9_inst_0_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_0_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_1_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_1_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_2_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_2_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_3_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_3_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_4_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_4_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_5_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_5_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_6_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_6_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_7_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_7_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_8_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_8_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_9_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_9_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_10_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_10_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_11_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_11_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_12_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_12_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_13_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_13_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_14_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_14_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_15_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_15_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_16_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_16_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_17_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_17_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_18_dout_w: std_logic_vector(17 downto 0);
    signal promx9_inst_18_dout: std_logic_vector(17 downto 0);
    signal dff_q_0: std_logic;
    signal dff_q_1: std_logic;
    signal dff_q_2: std_logic;
    signal dff_q_3: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_11: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_13: std_logic;
    signal mux_o_14: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_31: std_logic;
    signal mux_o_32: std_logic;
    signal mux_o_33: std_logic;
    signal mux_o_34: std_logic;
    signal mux_o_35: std_logic;
    signal mux_o_36: std_logic;
    signal mux_o_37: std_logic;
    signal mux_o_39: std_logic;
    signal mux_o_52: std_logic;
    signal mux_o_53: std_logic;
    signal mux_o_54: std_logic;
    signal mux_o_55: std_logic;
    signal mux_o_56: std_logic;
    signal mux_o_57: std_logic;
    signal mux_o_58: std_logic;
    signal mux_o_60: std_logic;
    signal mux_o_73: std_logic;
    signal mux_o_74: std_logic;
    signal mux_o_75: std_logic;
    signal mux_o_76: std_logic;
    signal mux_o_77: std_logic;
    signal mux_o_78: std_logic;
    signal mux_o_79: std_logic;
    signal mux_o_81: std_logic;
    signal mux_o_94: std_logic;
    signal mux_o_95: std_logic;
    signal mux_o_96: std_logic;
    signal mux_o_97: std_logic;
    signal mux_o_98: std_logic;
    signal mux_o_99: std_logic;
    signal mux_o_100: std_logic;
    signal mux_o_102: std_logic;
    signal mux_o_115: std_logic;
    signal mux_o_116: std_logic;
    signal mux_o_117: std_logic;
    signal mux_o_118: std_logic;
    signal mux_o_119: std_logic;
    signal mux_o_120: std_logic;
    signal mux_o_121: std_logic;
    signal mux_o_123: std_logic;
    signal mux_o_136: std_logic;
    signal mux_o_137: std_logic;
    signal mux_o_138: std_logic;
    signal mux_o_139: std_logic;
    signal mux_o_140: std_logic;
    signal mux_o_141: std_logic;
    signal mux_o_142: std_logic;
    signal mux_o_144: std_logic;
    signal mux_o_157: std_logic;
    signal mux_o_158: std_logic;
    signal mux_o_159: std_logic;
    signal mux_o_160: std_logic;
    signal mux_o_161: std_logic;
    signal mux_o_162: std_logic;
    signal mux_o_163: std_logic;
    signal mux_o_165: std_logic;
    signal mux_o_178: std_logic;
    signal mux_o_179: std_logic;
    signal mux_o_180: std_logic;
    signal mux_o_181: std_logic;
    signal mux_o_182: std_logic;
    signal mux_o_183: std_logic;
    signal mux_o_184: std_logic;
    signal mux_o_186: std_logic;
    signal mux_o_199: std_logic;
    signal mux_o_200: std_logic;
    signal mux_o_201: std_logic;
    signal mux_o_202: std_logic;
    signal mux_o_203: std_logic;
    signal mux_o_204: std_logic;
    signal mux_o_205: std_logic;
    signal mux_o_207: std_logic;
    signal mux_o_220: std_logic;
    signal mux_o_221: std_logic;
    signal mux_o_222: std_logic;
    signal mux_o_223: std_logic;
    signal mux_o_224: std_logic;
    signal mux_o_225: std_logic;
    signal mux_o_226: std_logic;
    signal mux_o_228: std_logic;
    signal mux_o_241: std_logic;
    signal mux_o_242: std_logic;
    signal mux_o_243: std_logic;
    signal mux_o_244: std_logic;
    signal mux_o_245: std_logic;
    signal mux_o_246: std_logic;
    signal mux_o_247: std_logic;
    signal mux_o_249: std_logic;
    signal mux_o_262: std_logic;
    signal mux_o_263: std_logic;
    signal mux_o_264: std_logic;
    signal mux_o_265: std_logic;
    signal mux_o_266: std_logic;
    signal mux_o_267: std_logic;
    signal mux_o_268: std_logic;
    signal mux_o_270: std_logic;
    signal mux_o_283: std_logic;
    signal mux_o_284: std_logic;
    signal mux_o_285: std_logic;
    signal mux_o_286: std_logic;
    signal mux_o_287: std_logic;
    signal mux_o_288: std_logic;
    signal mux_o_289: std_logic;
    signal mux_o_291: std_logic;
    signal mux_o_304: std_logic;
    signal mux_o_305: std_logic;
    signal mux_o_306: std_logic;
    signal mux_o_307: std_logic;
    signal mux_o_308: std_logic;
    signal mux_o_309: std_logic;
    signal mux_o_310: std_logic;
    signal mux_o_312: std_logic;
    signal mux_o_325: std_logic;
    signal mux_o_326: std_logic;
    signal mux_o_327: std_logic;
    signal mux_o_328: std_logic;
    signal mux_o_329: std_logic;
    signal mux_o_330: std_logic;
    signal mux_o_331: std_logic;
    signal mux_o_333: std_logic;
    signal mux_o_346: std_logic;
    signal mux_o_347: std_logic;
    signal mux_o_348: std_logic;
    signal mux_o_349: std_logic;
    signal mux_o_350: std_logic;
    signal mux_o_351: std_logic;
    signal mux_o_352: std_logic;
    signal mux_o_354: std_logic;
    signal mux_o_367: std_logic;
    signal mux_o_368: std_logic;
    signal mux_o_369: std_logic;
    signal mux_o_370: std_logic;
    signal mux_o_371: std_logic;
    signal mux_o_372: std_logic;
    signal mux_o_373: std_logic;
    signal mux_o_375: std_logic;
    signal gw_gnd: std_logic;
    signal promx9_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_0_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_1_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_2_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_3_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_4_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_4_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_5_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_5_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_6_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_6_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_7_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_7_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_8_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_8_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_9_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_9_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_10_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_10_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_11_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_11_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_12_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_12_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_13_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_13_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_14_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_14_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_15_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_15_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_16_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_16_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_17_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_17_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_18_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_18_DO_o: std_logic_vector(35 downto 0);

    -- component declaration
    component LUT4
        generic (
            INIT: in bit_vector := X"0000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic
        );
    end component;

    -- component declaration
    component LUT2
        generic (
            INIT: in bit_vector := X"0"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic
        );
    end component;

    -- component declaration
    component LUT5
        generic (
            INIT: in bit_vector := X"00000000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic;
            I4: in std_logic
        );
    end component;

    --component declaration
    component pROMX9
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(35 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_gnd <= '0';

    promx9_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_0_dout(8 downto 0) <= promx9_inst_0_DO_o(8 downto 0) ;
    promx9_inst_0_dout_w(26 downto 0) <= promx9_inst_0_DO_o(35 downto 9) ;
    promx9_inst_1_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_1_dout(8 downto 0) <= promx9_inst_1_DO_o(8 downto 0) ;
    promx9_inst_1_dout_w(26 downto 0) <= promx9_inst_1_DO_o(35 downto 9) ;
    promx9_inst_2_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_2_dout(8 downto 0) <= promx9_inst_2_DO_o(8 downto 0) ;
    promx9_inst_2_dout_w(26 downto 0) <= promx9_inst_2_DO_o(35 downto 9) ;
    promx9_inst_3_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_3_dout(8 downto 0) <= promx9_inst_3_DO_o(8 downto 0) ;
    promx9_inst_3_dout_w(26 downto 0) <= promx9_inst_3_DO_o(35 downto 9) ;
    promx9_inst_4_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_4_dout(8 downto 0) <= promx9_inst_4_DO_o(8 downto 0) ;
    promx9_inst_4_dout_w(26 downto 0) <= promx9_inst_4_DO_o(35 downto 9) ;
    promx9_inst_5_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_5_dout(8 downto 0) <= promx9_inst_5_DO_o(8 downto 0) ;
    promx9_inst_5_dout_w(26 downto 0) <= promx9_inst_5_DO_o(35 downto 9) ;
    promx9_inst_6_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_6_dout(8 downto 0) <= promx9_inst_6_DO_o(8 downto 0) ;
    promx9_inst_6_dout_w(26 downto 0) <= promx9_inst_6_DO_o(35 downto 9) ;
    promx9_inst_7_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_7_dout(8 downto 0) <= promx9_inst_7_DO_o(8 downto 0) ;
    promx9_inst_7_dout_w(26 downto 0) <= promx9_inst_7_DO_o(35 downto 9) ;
    promx9_inst_8_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_8_dout(17 downto 9) <= promx9_inst_8_DO_o(8 downto 0) ;
    promx9_inst_8_dout_w(26 downto 0) <= promx9_inst_8_DO_o(35 downto 9) ;
    promx9_inst_9_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_9_dout(17 downto 9) <= promx9_inst_9_DO_o(8 downto 0) ;
    promx9_inst_9_dout_w(26 downto 0) <= promx9_inst_9_DO_o(35 downto 9) ;
    promx9_inst_10_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_10_dout(17 downto 9) <= promx9_inst_10_DO_o(8 downto 0) ;
    promx9_inst_10_dout_w(26 downto 0) <= promx9_inst_10_DO_o(35 downto 9) ;
    promx9_inst_11_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_11_dout(17 downto 9) <= promx9_inst_11_DO_o(8 downto 0) ;
    promx9_inst_11_dout_w(26 downto 0) <= promx9_inst_11_DO_o(35 downto 9) ;
    promx9_inst_12_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_12_dout(17 downto 9) <= promx9_inst_12_DO_o(8 downto 0) ;
    promx9_inst_12_dout_w(26 downto 0) <= promx9_inst_12_DO_o(35 downto 9) ;
    promx9_inst_13_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_13_dout(17 downto 9) <= promx9_inst_13_DO_o(8 downto 0) ;
    promx9_inst_13_dout_w(26 downto 0) <= promx9_inst_13_DO_o(35 downto 9) ;
    promx9_inst_14_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_14_dout(17 downto 9) <= promx9_inst_14_DO_o(8 downto 0) ;
    promx9_inst_14_dout_w(26 downto 0) <= promx9_inst_14_DO_o(35 downto 9) ;
    promx9_inst_15_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_15_dout(17 downto 9) <= promx9_inst_15_DO_o(8 downto 0) ;
    promx9_inst_15_dout_w(26 downto 0) <= promx9_inst_15_DO_o(35 downto 9) ;
    promx9_inst_16_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_16_dout(8 downto 0) <= promx9_inst_16_DO_o(8 downto 0) ;
    promx9_inst_16_dout_w(26 downto 0) <= promx9_inst_16_DO_o(35 downto 9) ;
    promx9_inst_17_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_17_dout(17 downto 9) <= promx9_inst_17_DO_o(8 downto 0) ;
    promx9_inst_17_dout_w(26 downto 0) <= promx9_inst_17_DO_o(35 downto 9) ;
    promx9_inst_18_AD_i <= ad(9 downto 0) & gw_gnd & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_18_dout(17 downto 0) <= promx9_inst_18_DO_o(17 downto 0) ;
    promx9_inst_18_dout_w(17 downto 0) <= promx9_inst_18_DO_o(35 downto 18) ;
    lut_inst_0 : LUT4
        generic map (
            INIT => X"0001"
        )
        port map (
            F => lut_f_0,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_1 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_1,
            I0 => ce,
            I1 => lut_f_0
        );

    lut_inst_2 : LUT4
        generic map (
            INIT => X"0002"
        )
        port map (
            F => lut_f_2,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_3 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_3,
            I0 => ce,
            I1 => lut_f_2
        );

    lut_inst_4 : LUT4
        generic map (
            INIT => X"0004"
        )
        port map (
            F => lut_f_4,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_5 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_5,
            I0 => ce,
            I1 => lut_f_4
        );

    lut_inst_6 : LUT4
        generic map (
            INIT => X"0008"
        )
        port map (
            F => lut_f_6,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_7 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_7,
            I0 => ce,
            I1 => lut_f_6
        );

    lut_inst_8 : LUT4
        generic map (
            INIT => X"0010"
        )
        port map (
            F => lut_f_8,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_9 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_9,
            I0 => ce,
            I1 => lut_f_8
        );

    lut_inst_10 : LUT4
        generic map (
            INIT => X"0020"
        )
        port map (
            F => lut_f_10,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_11 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_11,
            I0 => ce,
            I1 => lut_f_10
        );

    lut_inst_12 : LUT4
        generic map (
            INIT => X"0040"
        )
        port map (
            F => lut_f_12,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_13 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_13,
            I0 => ce,
            I1 => lut_f_12
        );

    lut_inst_14 : LUT4
        generic map (
            INIT => X"0080"
        )
        port map (
            F => lut_f_14,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_15 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_15,
            I0 => ce,
            I1 => lut_f_14
        );

    lut_inst_16 : LUT4
        generic map (
            INIT => X"0100"
        )
        port map (
            F => lut_f_16,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_17 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_17,
            I0 => ce,
            I1 => lut_f_16
        );

    lut_inst_18 : LUT5
        generic map (
            INIT => X"00040000"
        )
        port map (
            F => lut_f_18,
            I0 => ad(10),
            I1 => ad(11),
            I2 => ad(12),
            I3 => ad(13),
            I4 => ad(14)
        );

    lut_inst_19 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_19,
            I0 => ce,
            I1 => lut_f_18
        );

    promx9_inst_0: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"E361B8E0703F180E880381D14C985C2D954B85A2892080412492072482194894522A190C",
            INIT_RAM_01 => X"E3E1F0DC804B2E16CA247228DC7453291408C3D1B0E0844B299449E3D1B0D45E37180FC6",
            INIT_RAM_02 => X"964B5D7E63077337598C461B0DACE87FBD9CAD25C2BD34AA54A812C7C34988C664359649",
            INIT_RAM_03 => X"45225974D65C3218CBF289BCC26F309CD26A551A954AB357A34E29349A853A7F42AA58EB",
            INIT_RAM_04 => X"E371B8D85E3121104844920128A45124928A4522914492482012080412410082412594CA",
            INIT_RAM_05 => X"C7B30944B45D319649E3E1F0FC704A2A16CA0461E8B8724A2893C7C3E1F0FC70411C1007",
            INIT_RAM_06 => X"148A7D165D38A556AA55BB1D82870877375A8C258AA974C46AB7196C15829D3E99542611",
            INIT_RAM_07 => X"E382092494492010CBA6C31970C65530A0B6B369C526A559A7CFE8140A4D46A34FA2CFA7",
            INIT_RAM_08 => X"E36178C06039208E882412090492422A148A452291249248201049248201008E38201208",
            INIT_RAM_09 => X"2B64EA311E984CA7D186A2F920945D321849E3E1B8FC704A299689E3E1A8D86E301F8FC6",
            INIT_RAM_0A => X"D3FA0522914E9ACD66F47A74F2492FA05227F41A954277087BB95A6BA58AA154BB663519",
            INIT_RAM_0B => X"04020924924124124945020104944A29148A4532A165089139DAF0D3FA052AB551A74DA6",
            INIT_RAM_0C => X"E371F0BC6E37180DC60381C8E8864B2994CA652249289241249208040201008041241008",
            INIT_RAM_0D => X"CD35CAA152B46AB79A4BE499ECFE914D29D1A712F93C8454321648C3E1B91C7E42259649",
            INIT_RAM_0E => X"D3FA054AB550A2CB24B36A0522914596C965F47A2CCA371C92CB64B269851E6712803C1E",
            INIT_RAM_0F => X"C371F8E08E38201048249249208E412492084522812494542C92CBA67502A55059B3E6F9",
            INIT_RAM_10 => X"C361B8E07E381D1206E371B8BC603921124944925148A452289208041200E08040238F87",
            INIT_RAM_11 => X"716945027B2384BE5F0F464AA14EAC6B39DC6BE4A211009A5527CF86A2C13C7243291448",
            INIT_RAM_12 => X"0A255AE1456CC6F5FFD3FA0D4AB550A2C8E37259FD02AF46974B65D35964AA230B8DC4A1",
            INIT_RAM_13 => X"0402010070471C1008040238E080471F8E08040201049048201008E4020928985A43A952",
            INIT_RAM_14 => X"4612B9187E39209207E361B8DC70391C904724120900824A2914492412010080402011C7",
            INIT_RAM_15 => X"9249144603088140A071594D0EA13C8D425F0FE71AD92C9B67BA5DAC74D9F1009A51278F",
            INIT_RAM_16 => X"24021940E2B257A696AC768CCEFD9DEBFFFFD3FA0D4AB551A6CAA251C9B4FA8D349246E3",
            INIT_RAM_17 => X"E382011C70471C11C7E382011C704124104924F1F8E08040238E080471F8E08041281008",
            INIT_RAM_18 => X"ACD449ACEC8047A10D451278FC6E312090070392090472412092492492490080401C0E07",
            INIT_RAM_19 => X"10B924B66D348D42A15098041DE10285C32271490D2EA75698C3DE3017F3614A9360385D",
            INIT_RAM_1A => X"E3F1F8FC7C37201048C6E4C26140A546A2D6CCCC0D972DEEFB7DFEF47A0D46A350A24AA1",
            INIT_RAM_1B => X"0402010080402011C7E3F1C10080471F8F86E3F1F8FC7C3F239187C3F1F8E08E3F1F8FC7",
            INIT_RAM_1C => X"51384BC9588856B3DA8B53D18CC8763B9F0C652249048242251249249249249249209248",
            INIT_RAM_1D => X"D3FA3D02934FA2486110081C765B2C8CC1DEEF77BBDDE30D97CDE6B249050EB75F98C3DF",
            INIT_RAM_1E => X"E3F201008040201008E381F91C7E42249E54E9852A310E9A57A8137B5C365FFFFFFFFDFE",
            INIT_RAM_1F => X"2492492080401C0E07E3F1C0E080402010480461B8E08E381F8FC6C371F8FC7E3F1F0F87",
            INIT_RAM_20 => X"D2B8F4C6A345903D9C0F27FB694E8F4A2D986A8471FD008A4823CFA6B2D148944A25148A",
            INIT_RAM_21 => X"989DBFDBEFF7FFFDFFB359B4FE8F3E9A461FAE6754565D3490C19E0F9833DDE511A1D4A9",
            INIT_RAM_22 => X"2381F8E07038238F86C3F1F8E08E3F1F8E070401F1910A804FA5D3A8D44AA962AF522330",
            INIT_RAM_23 => X"A722D14892492490080402010070381F8FC7E47238FC7E38238E080471F8FC7E3F1C0C48",
            INIT_RAM_24 => X"3018441DE712A6D92AD2A86C7E533F92C29E6FB823FDA8BD5FB21AED6622D166AB54A410",
            INIT_RAM_25 => X"E98512D922A934D930BD7FBFDFEFF7FFFFFE72496CDE7F3E96C61E8D57143E714694C01F",
            INIT_RAM_26 => X"0401C8E48238188F088491C0C4723A208EC8853280FC7E3E1B8ECA06D4AA013C9442A055",
            INIT_RAM_27 => X"2EF6EB3188B253A30E459241008040238E080471F8E0803F1F91C7E381F8FC7C3F1F8FC7",
            INIT_RAM_28 => X"EF07DC7E83409E441F51389439E3089950A8F2C8BC8A7B55A5D066331984BA390B7DBEDF",
            INIT_RAM_29 => X"A9546A150C90502951E9853A9D3D10B367BDDF7FBFDFEFF7FBFEF9314934C28349A04EE2",
            INIT_RAM_2A => X"C3F1C11C7E3F1F900703B21A05D121B8DC2C162BCDA6D36E8CBC15E6425908884A3BA592",
            INIT_RAM_2B => X"953A55026D2485C01EEE5612C55E963D988A2482011C7E3F230F86C3E1F91C8E3F1F0FC7",
            INIT_RAM_2C => X"51698D2AA54BA953E671181C9E71479EC86050B89C05E4FF91D16B955AAD7ED168BBDB6B",
            INIT_RAM_2D => X"D5FB14F9C0321E940D87E4B25D2C8E4E2111EA5482BF497FCFFFFFFF7FBFFFFDFEF6DE31",
            INIT_RAM_2E => X"C3E1F0F87C3F1B8FC7C361B8FC7E381C0DD4949B8DC6E578B7D82EF66AC5A2E168B45BEC",
            INIT_RAM_2F => X"381C0607037EB254A913E9644A00F772B2962A74FA34F86A2C964904F238FC7C3E1F0D87",
            INIT_RAM_30 => X"FF7FF7FFDF98CDAED7720A154AA554AE56A9B2984C324F3796C4E07058F47E4134ABD82E",
            INIT_RAM_31 => X"9529D50E974CAA55ABD5EAF562DD5A9AA70A03737251067C451F52A8B3CEB711A7FFFFFE",
            INIT_RAM_32 => X"040238E080471F0FC7E3F1F8FC7E3F1F8FC7C361B0D86E31385A6E165AED56A953A652E8",
            INIT_RAM_33 => X"73CAA556BD6FB8E0B1591C3DD6C5519F492350F7AB7196C25BA9D3C853E1ACC459281208",
            INIT_RAM_34 => X"433BEE2F9FF7FB7DFEFFFFC672F32E6A30D7929A658EB553ADD467D23854122F2898CA66",
            INIT_RAM_35 => X"953A252A7542A1D2A853A9CCEE9F67B2D6E953AA1532AD67B7D82D0EF3317CC68139A0D0",
            INIT_RAM_36 => X"A7B35184A248241008E471F8FC7E3F1F8FC7E3F230F87C361B0D87C371F8C060E8BBD96A",
            INIT_RAM_37 => X"338984C68954AAD7ACD6FBFDFEF17FBFDFAED75B5D6A9F348DC25F0F56DB0560A84FA590",
            INIT_RAM_38 => X"F629FAB43C662DA08F375C779FEFF6FBFFFEBDEC8E8556BF502A15D31A1D4AA343A654E9",
            INIT_RAM_39 => X"E3F180CA716DAE52E85499D4EA7543A550E9542A1506733A9D4EA853BA54E6733A9DD36B",
            INIT_RAM_3A => X"EF5692E150A74F230F66A2C944904F238FC7E471F8FC7E3F1F9187C361B0D87E3F1F8FC7",
            INIT_RAM_3B => X"13CAB59ACD5EB3DBEDD5DB2D9ADF77BC5FEF181C35F6E96BAD54AA552A8D228B2B8D425F",
            INIT_RAM_3C => X"5419C4E27F3797CDE533D88AC8E64222D2ADD9EFBFDFEDF7FB79F27BD4CAD9388D4F2793",
            INIT_RAM_3D => X"C361F8F86E3F238FC70381E522DB53A4CEA73329D50A9542A14EA753A9CCC6733A9D50A7",
            INIT_RAM_3E => X"D3FA3D1E7B248D401FCEC64ADD3C95421C8C4592412080471F8F87C3F1F0F87C3F1F8FC7",
            INIT_RAM_3F => X"02C411CD0A94472952D60B8DE6F379C16070180C06231D87C35F6E973B1D8AB357A34FA6"
        )
        port map (
            DO => promx9_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => promx9_inst_0_AD_i
        );

    promx9_inst_1: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F62A357ED7499D50683419C4C26F3696475C6842B960DE63BA60B7DF7FB7DFEDFFCD5C5F",
            INIT_RAM_01 => X"C3F1F0FC7E3F238F86E381C0C070301C0E4724344DB6A54198CCA8952A2552A543A1D267",
            INIT_RAM_02 => X"150A45229F459A48E491C92CB66B22843D5B6CA5FA750873349449040238FC8E471F8F86",
            INIT_RAM_03 => X"FF6FBFD3977BBDC1A22AC25918B6411C9C8F382C9E6F2592C966B2390C7E1AFB73B5566A",
            INIT_RAM_04 => X"5429CCEA73399CCE263399C4E67339A0CC271309FCBA530469210A64C26944ED4CC3F9BF",
            INIT_RAM_05 => X"E472391C8E472391C8C3F238E07E301C0E4844E339A0DE662C1AD00AEAA54A813198CE66",
            INIT_RAM_06 => X"D7DBE5CEC558ABD1A7B3496CB6592A88C21FEF285C7249187EB696E9C419A8C250241008",
            INIT_RAM_07 => X"8552846AEB8EF3FDFEFF7FBE531B56AF542D16FB3D82D780549D8B79ACD66B2188C3DFAF",
            INIT_RAM_08 => X"D56AED4E91319CCE6733AA150673409CCE673399C4C67130984DE6D2C8CBE9807526134A",
            INIT_RAM_09 => X"6692812090402391C8E47239008E47238E070432B180E8915C3B6333CA9D2E9954A950A7",
            INIT_RAM_0A => X"38FC75F6E762B1DAEC562AD566A14E9E4AE33007FBE1FEFE72B4D86C56FBC5F0F66DAD91",
            INIT_RAM_0B => X"EF05C1B4AA552B17CCC5AB55CB7FFFFB7BBE3AAB5D0A733A9DD0A874BA5512A746B3576A",
            INIT_RAM_0C => X"795D7F039DADAD50A974EAE61ADB64AD50A73399C4E671399C4C26F379BCDE5D2692C8E1",
            INIT_RAM_0D => X"A8744AB178C257A4CD2502011C8E47238FC8C3E1F0FC6E3B2B9D126C17C4B6AD5DAB57EE",
            INIT_RAM_0E => X"33AA1D2A9543A253ACB74B5D66A349A8542A157A34FA6B338CC1DEAD3652E572A8532350",
            INIT_RAM_0F => X"F2E974B6471286B9D50762F17CC06835A0CF364C6F5FEFF7FAF8EFD519CCFE6F2898CCA8",
            INIT_RAM_10 => X"F68B9E5B51C1E4F3F7BABC8DFECB509B49E4F2AA1D42FD68BF5AA93419CCE671309BCBE6",
            INIT_RAM_11 => X"09E469F0E873311449251259B4FC84391608E47239187E3F1F0FC6E381D944F0A978CD6A",
            INIT_RAM_12 => X"338984DA5F31A0CE6753AA152A874CA5D2E975AACD5E8D3FA3D1A7D3D9ACB245107A3296",
            INIT_RAM_13 => X"751A04E26F3797CDA5B258D4261ADD4F994AC5F33988FA9C64382B19EFBFDFEDF6CDE067",
            INIT_RAM_14 => X"C5E513F28D58BA66375D2E8F3B5789C05DADD66B2D8EA1379749A4F2898CF2B179C1636C",
            INIT_RAM_15 => X"D3E9B4B232FD6BA70E66229148A24924924904928944A2482791C7C3E1F0FC7E371F8E07",
            INIT_RAM_16 => X"FF6FBFE34778944D6A3319CCFE63399CCEA7543A550A954BA5D2E9140A3D1E7D369B4DA7",
            INIT_RAM_17 => X"F2F984CA8178BDE333D6AA04E26F2E96C923711823552E652A134AC5F3223D46CFAA5EF8",
            INIT_RAM_18 => X"4532A97CD075301C5690DA85B743B9E06FF6999C05DEDB65B2D96CD68BCE1ADD63A7C9A3",
            INIT_RAM_19 => X"140A3CFA6D369ACDE7F3F9F4AE2EEA5A9E4A249249249250241208048201249249249249",
            INIT_RAM_1A => X"E623EA511D46CBFBFEFF4ED5BEB9158BC963D28984C27342A15067542A150A854BA5D32A",
            INIT_RAM_1B => X"182CA69B6FBDD15163B2693CC67D6AE3ECB1183A84FE5D2D92441E6CC47994A84C26958B",
            INIT_RAM_1C => X"65E3820916944F29D62C36632970AD6BC76B37FD4F1F5992BC5FADD6EBB5D6DD6FBC5E70",
            INIT_RAM_1D => X"339A152E954BA5512A140A34FA6D369B4DE7140A3CD23EE9559849248201009048201048",
            INIT_RAM_1E => X"C6426130984C2A954A06C4231691AFFFFDFE98BBF36A070D8F4764D2797CBE5F309C4E68",
            INIT_RAM_1F => X"D6FBBDFEFF78B85FEFF70BCE2F3FC1EB6C26B258F4A2674BD176FC1C8C0D027B217DB311",
            INIT_RAM_20 => X"2482494CBA67349F13EB36AB9DE2FA8647A4F2E943D9B90DA961F61BDC8DBECD65B2D96C",
            INIT_RAM_21 => X"B1E934A261319C4DE51399D50A7542A1D2E9147A3D1E8F3F9FCFE8140A34CE2CDF491608",
            INIT_RAM_22 => X"DFCF0D364AE6541B0984B22130984D281A4EE5F8CDCB7DF7FD6CEF6FE6FBA1E50381C321",
            INIT_RAM_23 => X"F65A9D32B965B2DB6C964B1D72C550A3CFA6D369850AAF7FE2FBADD248EC9A5345D77DFE",
            INIT_RAM_24 => X"348A04EE1CD9531D8D07A4227952C36C3EA1B2798D0A9553A5D52B75490BEE7176D46EF1",
            INIT_RAM_25 => X"0A959B15AEE17941229148A4563D279749A433898CE263399D50A8148A051E7140A05028",
            INIT_RAM_26 => X"91C89C563D2AA7FF3CFFEFBDED82742590C864321914A072411F10731D77DFEDECC5E152",
            INIT_RAM_27 => X"71486D5321BDCC5929542A257ADB64B1D6AA34698C31B0B4491E4F47B46A6168D07EC9A5",
            INIT_RAM_28 => X"349A45028349A4D069349A0CD618F1682E988DF74C0E2B20A1552CB6DB75DEEF77BB5AEA",
            INIT_RAM_29 => X"7C7FFFDF4D5031A111A97512ED98D673BA5F50485C0E070D8A4563D2690CE661309CCE67",
            INIT_RAM_2A => X"84C26134AC58392153EAA62379E71697EF76192CFD108643210E8743D2C1CD168F36BE6C",
            INIT_RAM_2B => X"181C06030187BE56A0D1FB76BF636EA9D2A954AA6572C552A851648DC4F170984C261309",
            INIT_RAM_2C => X"50384BEE1917944A67552A954AA341A0D068544A751A6B248E47A5132A1D56CD77BC5E30",
            INIT_RAM_2D => X"E734624D1C6193653AFF9D55C65C5830188EA8C47ABD56C46B39DD2F97CBC5E5017CC05F",
            INIT_RAM_2E => X"A542590884422110874421D10876432190C864D2F184F68A41A313E6C2590874421D10C9",
            INIT_RAM_2F => X"F78C0E2B1592C964B258AC4E270184B1C3E4580DF686CD53A5D4A974CAED8EC34D96BB12",
            INIT_RAM_30 => X"EE673375B6CB64AE970B05BAA164BE6CBD63752A954A9549A05067940A9D76BB65B2D9AD",
            INIT_RAM_31 => X"6421C8E462311A149089551A2D7118CFFF7BD99958FCBC572F97CB2723EA5940AB62335B",
            INIT_RAM_32 => X"B67C0E5F09205F9AC96421D0E47231188C462311C8C46231180A46231188C062321D90C8",
            INIT_RAM_33 => X"941AFDEB158AC562B1794CE66F379AC96472592C4E23096488CD321C5CFD76A953A9D52A",
            INIT_RAM_34 => X"0623D2153A9A5D2F194C15B291188B3D1E4E2693419CBC572C1752752A4D268340A04E26",
            INIT_RAM_35 => X"028140A05028148C46230180A052352DA3138903A3E6E9C7FEE3612AF2E954AE5D2717CB",
            INIT_RAM_36 => X"987AF556A954AA57F059ACA5AA2AA4291047231188C05028178A05028140A05E28178805",
            INIT_RAM_37 => X"349A050271309BCDE5943B463349A4D269339A4D268F3591C46070389C4E2EC90AA2E877",
            INIT_RAM_38 => X"A552A930984C221109A4F2DA111895482A56EAC441D8BA54269349845269349C4E2B13CA",
            INIT_RAM_39 => X"C26130984C26130BC4E271389C4C27138A05E2F138BC56493DA2D288F8BE7BE3AEA7A78A",
            INIT_RAM_3A => X"178C2D963336D06CF0F5FAF552A95DB3DEB259CB3BC90852208E460281789C4C26130984",
            INIT_RAM_3B => X"83C1E9149A4D269349549A4D06713F9BCBE473AB0E334BADD6693379BCDE6B217EBB5BEE",
            INIT_RAM_3C => X"36BE3FD710A62B974AC562A954984B2210C88462C1A8F88D4B27946803692C763B1E1107",
            INIT_RAM_3D => X"E271389C4C260F0784A1D0E8743A1D0E8743C1E138984A1D0F09C4E2F138805E67591FDB",
            INIT_RAM_3E => X"79BCD6471B62A4CEA8962AB48A7990DAE570778B357ACD60C26AF496E74A0C94411C8C05",
            INIT_RAM_3F => X"E6C258EC763B1D8EC763B1A0F0784526110895BA9D26833F9747A3732B0E574BADD66933"
        )
        port map (
            DO => promx9_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => promx9_inst_1_AD_i
        );

    promx9_inst_2: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"E27138A88EB1314BF2DDDE5BF8BC552B1549A5426130984421908743D26114A27B4222D1",
            INIT_RAM_01 => X"EF2469487230180BC4C260F0983A1D0B0743A150E8702A1D0E0502A150E8743A1E0F0984",
            INIT_RAM_02 => X"72AACE374BADD2E93379AC8E3AE34488BC5E2EA804CF13BECDDEEFB8BC0DCB058DDAED6E",
            INIT_RAM_03 => X"43526130884F349C4EC5C210C8663B1D0C8663B1D8EC7633198F07B64AED72A7499FC962",
            INIT_RAM_04 => X"A140A8743A150E8784E2F100A874ECB9F1FE9835B174A84C26114984D26938A84D299087",
            INIT_RAM_05 => X"984C6E532DBFE35E2089D2D104602F1789C4C1E0F0743C1D0E85028140A03018150A0302",
            INIT_RAM_06 => X"D6EB3596B9529FC961522A8E575BAED6E934791C75CA87066E30D8ACF9160371B5C66130",
            INIT_RAM_07 => X"84C221308A4C2292C843A190EC743A1F178B642188A4522A190C8622A190C86431148A86",
            INIT_RAM_08 => X"2360D82C080B0583018140605028150F0784C20149BA9967FE72A606036954943A1E1149",
            INIT_RAM_09 => X"916B2E635D9BBE6173DA6D2E9F8FC2D24995E6A208C46E27130983C1E0E05422352E9509",
            INIT_RAM_0A => X"228108A45021148A45F6FB357AB952A04760319A46374BADD6E8F3596B8CE5FAD461AED7",
            INIT_RAM_0B => X"E662E970884422130863B210EC784C22110984A198E46028158E4722914084522A188A45",
            INIT_RAM_0C => X"64C67442432A9449E3D0D813BD3A481500C060C0602C180C068784E2657D3BAFF7CA33CB",
            INIT_RAM_0D => X"D719CBAD86BA592E5EB54C46DB4784C767B4DA6D06F3D9A89D32908511C0C05E27130983",
            INIT_RAM_0E => X"228108A04228108A45220100845E20100805370B7D9ABB529BC51EF079F5EF49A3CD6430",
            INIT_RAM_0F => X"525EB7FFD16546134AE65299109644219108644208C4643426134A840140805021140845",
            INIT_RAM_10 => X"438178BC4C2713221BB047CB81B0DA753A9D6F072B318CD66AA3CA23201008160C068414",
            INIT_RAM_11 => X"8EC965A71186BAD8E913B85B0974BA5B34A778FD86BB3B98D86CF198ED470FC3957627CD",
            INIT_RAM_12 => X"C1F1389C40201008040201008040201008030181387C3E1F0F85C3371BBDBAB94092C09B",
            INIT_RAM_13 => X"C802D8FC4C143F4EB5BDFFFFC9EC52190F09A55299086232190EC76432283C363A1990C8",
            INIT_RAM_14 => X"1B1E06EB171F581EC90301789840A871BDDA0D86D3B1ED0F8740DD6B43B8D45A21089A94",
            INIT_RAM_15 => X"369B859AA73789BBD80C9844EEB7509AC72290C8A42E09117B462EDA7D6E572FA1DEE973",
            INIT_RAM_16 => X"43B238886A0A1F07C3C1E0F87C3E1F1386040201009C3E1F0C09C4E200C06C4A2A0E8542",
            INIT_RAM_17 => X"0401F0F86C351A0842476653A23158ACE738BCCC2A384E20150D8AA552A128743B218E87",
            INIT_RAM_18 => X"D9BBDDF71981BBEA783C0DC5D242C246968702F12A45D4F45FB21B6F57FC5E2D0271AACB",
            INIT_RAM_19 => X"C240B8A88037138B84368B3D7693247C3355CB36940261358D4162133AAD76B7499A5332",
            INIT_RAM_1A => X"6432190C822B1D8E864321D91C463A1A8583C1D0B0582C160F89C3E1F0F8404215120703",
            INIT_RAM_1B => X"8FC7CB7984A4378E08E3F1F0D86C36160A84216039316EDA97D46C73D2F0783E20140AC7",
            INIT_RAM_1C => X"D61C162F1D62A0DFB477EABD62B943C0F036BA4ADC51A89F35944643276C1166B567B21B",
            INIT_RAM_1D => X"C1F0F8883616160503A240E0744439198CC5360AC576931B732D1489F5B38A0B17944EA9",
            INIT_RAM_1E => X"E250A8583C1F100A0543B219087028150E05432190DC3010070302A150A8342C160F0783",
            INIT_RAM_1F => X"B0A75AD17CC86BB5174AD3D9A4AC361F8DC7C34178DC6A2A0D044200E0303C1A835AC01C",
            INIT_RAM_20 => X"696573922333AAD62F795CE64B1B5BA15EF0D54A057A9167D3E8B013287BC17686319192",
            INIT_RAM_21 => X"60D0A8341A150A8542C1D060985E240F0806E2E1307838431A0D88369B057A831A6EAAD2",
            INIT_RAM_22 => X"00D0281408033B254260C0A8502A1F1389C422A1D8E86020140A8743A1C8502A1E0E04C3",
            INIT_RAM_23 => X"7087E379527C2BB7A26B255AD58CCA561FC8C3E1F0D45A35168BCFEE584B714E69260B00",
            INIT_RAM_24 => X"772B4D96931A72AB554CF7AC62674DAC5C70794CE67EE333A45A2D53A99D02BB8CBFD7E5",
            INIT_RAM_25 => X"C0F030BC5E101282C140901830280C0685426050D8383E27138A46439180707C47228C49",
            INIT_RAM_26 => X"3329BC49DAAF3A1585E0B0302C04020290C1403018301A17138983E221D8E04228140A46",
            INIT_RAM_27 => X"53A9B55B256BA3C8A10FE753313E627B42534B562B09566D1988C44221209056271C3CA7",
            INIT_RAM_28 => X"A4D1F0F45E4719954B77BBD5C2B7357CB31A0FE91536BD66B35BEE58CCE656B336AC5B6A",
            INIT_RAM_29 => X"E21188C874391B8B00C04088A860191385418120100C060B0682C340B070983E20150D49",
            INIT_RAM_2A => X"41A0C86822407049A212580B61827E35944883C2901804030201014020102C1C1F130783",
            INIT_RAM_2B => X"58CCDE7AD536AF54E832C9E5FEC3358D405F0F5702ED2B057C24D56B45FA5CA4220D0883",
            INIT_RAM_2C => X"E260F888542A1B918624B299309E311E138A985C25EADF4A90401FD23A6D7ADF6FB45C70",
            INIT_RAM_2D => X"4020480C1A160F0783C18150E0502F1980C3A18150C844210C8602C0D0502C0603050704",
            INIT_RAM_2E => X"29B398A8341A0C864201007814CCC3753819EB967AF5427E2D9088C462603C0E03018141",
            INIT_RAM_2F => X"F2BA6D7EE382C562B299ED6676B32CA6502452FA5CFA391380BE1ECED6C2F608F1512916",
            INIT_RAM_30 => X"E150582004060C8D83C1B050B48C38259509644221348258311CD0B86C6E12F55E9ECB22",
            INIT_RAM_31 => X"6241908012050100802010080808160B0783C1E0F05C302B010502C1A158AC5423110844",
            INIT_RAM_32 => X"CEB67C55F29B55AA5446B1486832190803C1E0E0214D4AB65E2B54CA2409A8F26E2D9007",
            INIT_RAM_33 => X"D86C2E12D559A44E67544ABDCB19A4D2EB75DAED9E6EA53A994C6452996C3227097CBE1E",
            INIT_RAM_34 => X"423120D068310D8A43E16020040011110BC3E1C1892C96673B154A0672C968C4633A9F11",
            INIT_RAM_35 => X"06D2B168F27939914BE35258CC020702808060100808060D0B0542A0E0B0582200060604",
            INIT_RAM_36 => X"53589C3214FA7CBE1ECDF8EBE536AD5D2ACD82A0C86420100783C1C000720D3056309D10",
            INIT_RAM_37 => X"46237A213E984FA5D5B74B1D6AA554B2D9ACD6FB56334BADD6EB75BAED9E4E933095CD28",
            INIT_RAM_38 => X"805060340E050C88C482C168F068341588C501603814524E1888C52471F8ECA6423FA80C",
            INIT_RAM_39 => X"C0619AD17A7329984FC603624594D862ABCE84A36A340A0000010060100808060B020341",
            INIT_RAM_3A => X"DB6DCE2A8130954C65F2381C09F5027C3FDDB1680A6D5ABC56A187419048200E0E030180",
            INIT_RAM_3B => X"E31220647656301B948844026562B360ACDA961A3CC2654EB45E71589C5E534BA5D6EB75",
            INIT_RAM_3C => X"40000808060C020340A0C058082616090884834168D46A3D1A0AC3015030A47851211089",
            INIT_RAM_3D => X"2080401C0C06030140A061724D6E8F4114100783922D2AAE622B14A611F1041A04000000",
            INIT_RAM_3E => X"79BC9E6F399CD2EB75DB6D7DE6612E8EC5204FA7D3E9F4F97C3D21D05562997AB14E1B05",
            INIT_RAM_3F => X"215339F12074269447656170A47A57301AD06826B3B5DAD95C2C98756964563347B96533"
        )
        port map (
            DO => promx9_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_5,
            RESET => reset,
            AD => promx9_inst_2_AD_i
        );

    promx9_inst_3: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"E742B8EC1206060080A010080804030203418020D034380A118AC56251A8D46A3D1D8882",
            INIT_RAM_01 => X"4DD532D978A94894820000001C0C0603018080516208E434210B0D85D37B059A54241E91",
            INIT_RAM_02 => X"7569140E2135B060F379AC964F39A5D76BB6DADD75A25F22813E5E2F27D3E9F2F9783B60",
            INIT_RAM_03 => X"82C168D87C38260841C05301C0D2793F9B0B64A2192C8A48349AD106839A91D4DE74415C",
            INIT_RAM_04 => X"630231D4BE652B1491E642D1184410060080E0101008060406034161E0D8E020100C88C5",
            INIT_RAM_05 => X"2F1793E9F4F87AC11DAA75831D7AB14C1282208038180C06028140A0A0B144DC2A0902C5",
            INIT_RAM_06 => X"CAE35345ACB266BADC96099405F712A7DCB2592C562F299DD2EB75BABCEDBE5B1A7C3A5E",
            INIT_RAM_07 => X"81710080241D0508C4A34170F8804E220A42805351E9164C489E0EC67140CCA69346869A",
            INIT_RAM_08 => X"E05028487230010244A3B1F910B082401C906942593C6A190680C02000080C04040581C0",
            INIT_RAM_09 => X"390C155A390877BA1E2F178BC5E2FC86BFD6CA85CB019CBA4C9301A160A8542A0E0B8701",
            INIT_RAM_0A => X"E752F184FCB5559A542871C49CFEB5502E58B69A1C3DE3079ADA70589C06071793CDE4B2",
            INIT_RAM_0B => X"E000080804030107C0C1F0C04434220D06C4624168D88833110601C0049A410279439A0F",
            INIT_RAM_0C => X"C361A0AC5623150A02A0F038183E502E0703A102298556A845249005E2A1487C220B82C0",
            INIT_RAM_0D => X"186BB5BEE179C4E23118EB84F224FE73361D0E9783C1E0EF863B950B960B259EB33B91C7",
            INIT_RAM_0E => X"8020096102803B9DCDE6C2F9B8D0752A8AC0675058954AA8622995D6AA5C5DE0FE965830",
            INIT_RAM_0F => X"A4E2F990803B1382C0E00008080407018301A080906432190D0884833158AC56220F8340",
            INIT_RAM_10 => X"4CB6A3698E74251006E361B0D4582B1489C2C010280C1226260504A351A9E90EFE6E1C95",
            INIT_RAM_11 => X"9589D419CEEB88D36CB6CB2576DF78C0E23118DB44D625077339DD0E877BBDDD17832A17",
            INIT_RAM_12 => X"4231588422170681404010180CCC6C2E99CEA6736174B6142B994A62116014DCB040A0D3",
            INIT_RAM_13 => X"03947B0DCEC38E485FC7632968A04B170280601010080A0A0B0541E18110844422110884",
            INIT_RAM_14 => X"2F777B99BD04732858CE87C3ED5C531D908803F1B0D86A2C118801E13028180A0F080889",
            INIT_RAM_15 => X"42101810CABC4CA38E34E97BCDA8D9804F2CD6DB259ADF79C564F217F9A41A370978BC5E",
            INIT_RAM_16 => X"4281006432210C8602422108402E0E028100007000000057269ACB44B2592C985C291289",
            INIT_RAM_17 => X"E0D04014040E088B4CA3E3C18D247F28974DC822997464260901C02010080C1C0B068341",
            INIT_RAM_18 => X"D297E41637038243217027C3AE0AFD57AC99CE980BE92C542210882411C0FC7C3D158882",
            INIT_RAM_19 => X"E3A24908823A25948965100128A25A29160834E97BCD98D97C4F6CD77BB5A2F38BC963AC",
            INIT_RAM_1A => X"0020180C060D0409C38070B83C22210804024270781C1A03060180400008000004101186",
            INIT_RAM_1B => X"64B2512480461A0882E04000140C01060341C1D4E934C2D579B50FC53170180602038040",
            INIT_RAM_1C => X"389C05E2F386B8D09FEE381C25F2FA824322B14853FE2AF4502F1BEF07F364FE5E2A9509",
            INIT_RAM_1D => X"4010000000030289C6A1F1A8808E3F1F8E4703F080E0804E1F0CC234F983F1BAD980D1AE",
            INIT_RAM_1E => X"C220180802060000404020202C06060B0403C170785C1E0E038580E0E020140601010140",
            INIT_RAM_1F => X"EF076AE8F26F2C178AA542A14CA2461604810050181C0603028001203020543E281593C4",
            INIT_RAM_20 => X"75AA6C81EEEB84D1EE389C3DFAE9658F39DC0F17BB99CEE97D3F219148A42246DE54B11B",
            INIT_RAM_21 => X"A040180804050281C0E0B05810160B00800261B1106C461C120945A2C12890582B130380",
            INIT_RAM_22 => X"60402014000A0100402010001804000000402030286C2811028382A0D028181C0E028140",
            INIT_RAM_23 => X"70B87C823AAF59359D0F87EAB1147230980CC562E950A24F1A0482005018000801008080",
            INIT_RAM_24 => X"62315888400A018100752A6C81EEEA83CDAD389C6DA6830467B9DCCDD6F379C0E97D40E1",
            INIT_RAM_25 => X"81C1301008030200806030100408010080C0A160B84808060B05414060701C24190484C4",
            INIT_RAM_26 => X"E05018000A01008040404020140A06030180E060200800000081C42101E804A4581E8744",
            INIT_RAM_27 => X"AD66F381D0E874BE9F502804BE369F59B59D10779A91067130980BA4B21908A03E158640",
            INIT_RAM_28 => X"A0C058100A0212804221A10860020201014175AA6C61EEE97C4D6C180BC4DDD8CE6F375A",
            INIT_RAM_29 => X"C43020B42441188D84C240985C08020100404000000C0003028342E160B878280D078781",
            INIT_RAM_2A => X"642208E48E35150601C05010000A030500402020100806030582C0601018240002139186",
            INIT_RAM_2B => X"D6AA7BD5ACDD6AB55BCE773BBDDEE8743C1E2F07B472028E54B39D0FF7E295187130178A",
            INIT_RAM_2C => X"E05028382C0C0785828140180808010101C06040080806030582C0962A6C7DDCE27FCB2B",
            INIT_RAM_2D => X"8030001842491C8B82224060E8562B1C8A44E1F160481E00000000A05020000002060100",
            INIT_RAM_2E => X"310872F1046D27170A242209008C3D150801C040101C08010080402020100802020182C0",
            INIT_RAM_2F => X"F7BAF485F0EA7F486834282B59B8D56AB59CEE777B9DCEE777BA1D0EF76425D28D5533DE",
            INIT_RAM_30 => X"203030000E00018101A0B02014160C070741A0C060101802010080E000201002090283C0",
            INIT_RAM_31 => X"203038040401010040E0508958822C1E0D08608058B478351D8C8502712028040F0180C0",
            INIT_RAM_32 => X"EE66EC25DE845030DA8E4762B1107322954B4471B0B4582C118842C04008180801008040",
            INIT_RAM_33 => X"E000281C0E0D000242395B04EE12F27E47632F56B375AAD56B37DCEE773B9DCEE773B9DC",
            INIT_RAM_34 => X"0191704C1400030041204028180A07028040C0204808040301014160201808080B010281",
            INIT_RAM_35 => X"8030001C080100004080001010080402004320D3EB04EC3E218DC761F1A8D87A46231148",
            INIT_RAM_36 => X"CE66F379CCE66F399BCDD6EC25CA724AAA170C060A711E671910C923D1A8CC442A150B82",
            INIT_RAM_37 => X"406078280403008040A0E0405806060104C2596B8D1632F97D3E1ECD877375AAD66FB9DC",
            INIT_RAM_38 => X"242281208E3F1B11888301089C3809038040003020140806030000E00038100609008000",
            INIT_RAM_39 => X"E3C1609042200C89828030081C0A02048140604020040C060309C22351F0688E40291646",
            INIT_RAM_3A => X"2F772B75ACDF73B99BADD6EB79BCDE6EB79BCDE6EC29D86F3CA5148AC57A51106A299488",
            INIT_RAM_3B => X"0070381C0802028341A0F040282809008040A090F82020120C818459FB8D1642F9783C1D",
            INIT_RAM_3C => X"A191C8EC965431920784A211088239200DC7C3C190884E1C0401400040180C08060301C0",
            INIT_RAM_3D => X"49B4E24D106E3E9A48C3D150A44229100981A0B0081808010280C0E170702414150D8D45",
            INIT_RAM_3E => X"59EB951A44FF743A1D4FF72B55ACDF73B95BAD56AB55AADD6AB79BCDE6DC160E8D371E11",
            INIT_RAM_3F => X"20302808080D020100A040300808100B8340C050000C320F048140E090E0BC261E1289C5"
        )
        port map (
            DO => promx9_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_7,
            RESET => reset,
            AD => promx9_inst_3_AD_i
        );

    promx9_inst_4: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"C090A070441A138F0884B261689E662C2648C0C21910964B21104803F220A8501D050100",
            INIT_RAM_01 => X"AD56BBBE32EB2E1B8F089492210E6A2917C882A1007C2E1F0C0782A030081C0807038243",
            INIT_RAM_02 => X"E0D1907C3209180706397BDD5E570F703A5F2F56E335AEE773375AAD56AB51A8D46AB55A",
            INIT_RAM_03 => X"6471B0B052260901C04020200C0604028140A03048302A110003C281B090302612050500",
            INIT_RAM_04 => X"80A0001C0C07098945A290A0986C32231B8B6533C23CD4873DA24C4662A92C864C26150A",
            INIT_RAM_05 => X"8D46A35198CC6633198CB65B16290539994DA753B1D4FE70291BCA8290B034060C068340",
            INIT_RAM_06 => X"A271008C8C1C0982C0201028004E361C948938FBE542790E6CBC9FEE469B35AEE773375A",
            INIT_RAM_07 => X"E6236200DA4F2E9349642208F456270600006020180C06040200C200204098360C170680",
            INIT_RAM_08 => X"6270A02C00010581016020001808010E8DC8E3920900B84A4A261320341AB55EBD4D2154",
            INIT_RAM_09 => X"CDB61B15AEE66EB51A8D46633198CB61B0D84C361B19BB0A79148B45A2D940DC69299D8A",
            INIT_RAM_0A => X"0050E8742818188000C0B1E100422012808120102810782A2B9D8C186BA55E690E693CDF",
            INIT_RAM_0B => X"29D3731D7EB85F2C8723C42248F48733198A8442991C76180E8480603018100A020B80C1",
            INIT_RAM_0C => X"6532812CB6682397054180683416020180C0401038000E12120A080432A96CE2A052AB97",
            INIT_RAM_0D => X"F86BA562670E6D3EE0AD365B15ACDE6EB5198CB6632D96CB6130976C361B0972FE8E410D",
            INIT_RAM_0E => X"4020100002070100C160C010401C231F0589845228F8883C1D0A8640B08810324C2F9CD1",
            INIT_RAM_0F => X"24A249A138C052ADD76E788B6DE0C75CB02305A47AA11C2C459E8D05E2A9447C23128280",
            INIT_RAM_10 => X"6C36130970B27F44DECAF3411C784F2A8EC421107834080B0180802070280C0A090E8DC7",
            INIT_RAM_11 => X"837050784C003FB0D3F86B5D4267066DBEE0ADB61B119AD56AB5196CB65B0D94C25D2E98",
            INIT_RAM_12 => X"899341B0A44A090000402018000201008084C051084476141E0FC9C3E27120A057269148",
            INIT_RAM_13 => X"E070300C10100A0B4846334A0D56BD66AC1A0D1603058EB2903200CA75BADD60BC52A711",
            INIT_RAM_14 => X"6CB65B2D84C25D2E984C25D2E570A859B1DCCBE60A9C7E331E8A83000040380A04018080",
            INIT_RAM_15 => X"C1A2D9A8B25B338E0904D168B0A0824EAD60F7EB9D5E690E6DBEE0AD2612ED8AD56A3319",
            INIT_RAM_16 => X"2C95EB397ECF5B2F98CC452298DC7E0E0280402020080001008440C31241106A40269080",
            INIT_RAM_17 => X"20803010080B0180802070280C0E080D8BCB264339DD2EB4630852ECD5C309B2CF5CB54B",
            INIT_RAM_18 => X"AD15CAC988CC65B0D86C365B0984BA5CAE974BA5D2E560B057A912A925B25C68150D0882",
            INIT_RAM_19 => X"01B1F0540E4F2792CC66B0301D187B3E1CCC65826898C28556BFD7F85B553E59176DBF20",
            INIT_RAM_1A => X"0955A3B1D6DA683059F318E25B30ED64361ACBD552A54A17000080400018141E02148CC6",
            INIT_RAM_1B => X"47A321084A14038442217030140803008040006018080A0E088948262319A96EAB3C0A53",
            INIT_RAM_1C => X"F7DB5D42691770BD20CDA5C2A566C3612E974BA5CAE560A8582C972B95CAC16EAF56A6D1",
            INIT_RAM_1D => X"003018603A040F8A42E8F64A4CB253370ECC653529DD22AF4EA111A6B360D4B49E63B3DA",
            INIT_RAM_1E => X"0623B2794A9443A5488B563B1564D05EACAF91A5FAADEB12573255EC96C254300A010080",
            INIT_RAM_1F => X"0B0542BD5CA54E248F4772C11442110401C0E0F028100602008000E06020000A0506830A",
            INIT_RAM_20 => X"8612B9548C7663329DF86BA56A8D2077B8DF0EA5FA9D42B25CAC160A8582BD4CA653AA15",
            INIT_RAM_21 => X"ABE4C0100600010080262098844E291C018A01D4094CC46A2F8B50A7746B1D2E9C60ABD3",
            INIT_RAM_22 => X"0070281C080401810223D2E28DDEBE561FD3E514CA61A4A26E3E66F7AA3B5590FF95C399",
            INIT_RAM_23 => X"CA6532994A9E4F29D4EA6532993A9449A08FE6B2C8F8461A0481C0C050200C0402008040",
            INIT_RAM_24 => X"29848A8D72A84E1ECBC7D371D8126A2AB0D518EBAD8A9F317BB8E04FB632953EA0542B94",
            INIT_RAM_25 => X"2997FB6954AE5E9B5062E018140C04018080E3F1A088AA601F3C91E7C2E194DE86022548",
            INIT_RAM_26 => X"0170301408030180802000301804020080004101A185209A328F47A782D18CBA7542AF17",
            INIT_RAM_27 => X"4FD6BA912A964EA752A954AA753A9C4AA793C9D4EA51288B409F0E8762D8E45C1C0D0440",
            INIT_RAM_28 => X"C753714CAE5648BA548B459AC952AA52A20BA7A321480A042E2E16F86BADAEA13387B89F",
            INIT_RAM_29 => X"00F200F4602E101089E7D3497878471082C0A0700008120F030140819208C0343C27114D",
            INIT_RAM_2A => X"2783314C72350A0280208030180804018080200038180001008180002020384E41090780",
            INIT_RAM_2B => X"F85BA58EA13B8B381D4FF702B1188D4A231188C45A2D168B41A31189445A2D04793C9C4F",
            INIT_RAM_2C => X"43B1B1309C1B38A3972861E9C0646C5896D6ED6613CD56B747A1DAA7230040060C0700D7",
            INIT_RAM_2D => X"C02050040416038140604018000E30178742C13010083601000082E0C0A8542A1B0401C0",
            INIT_RAM_2E => X"482411E4F27034194F6793395482360E0281208030180A04018080401038180C070381C0",
            INIT_RAM_2F => X"C751F8080805030180F86BA56A912C8B379B0E875B11268341A0D068341A08F47A3D1E8F",
            INIT_RAM_30 => X"2221409C34360C01C0EA21E9989A8338268BE9D2E9652CBA4E9C5EED666B2566AA5014D4",
            INIT_RAM_31 => X"401038180A050301C0C050381C0C050281008040002402020081C0C04008080C030A05C4",
            INIT_RAM_32 => X"47A3D1E8F271389C4E47A3C9DCD06F3395CFA7B34978962F0A8682000038380A04018080",
            INIT_RAM_33 => X"0ED663014E9F4FA0958671C0100A0000804018FBE56A9F2C8BB99A0E97737D447A3D1E8F",
            INIT_RAM_34 => X"007010180006140884633150A804360A0281059140ECB47F2127DC92A2533614A48B2E8C",
            INIT_RAM_35 => X"00F0200C0803018040207038140802018140E06028140A030181000030182C1A13030000",
            INIT_RAM_36 => X"EE178BAD888A3D1E8F68341A0D047A3DA0D047A3C9C0D06E2C14500953D19CA4360D8240",
            INIT_RAM_37 => X"8AA5C3692AB9743399CCF6DB7990DB56AF0EE07220340E0D010302390C6D8A912D883B9A",
            INIT_RAM_38 => X"C0D0180C0A0D0180C1600018001810120C03833158A85631170500C392D2C96E6C54345C",
            INIT_RAM_39 => X"2A036820160B0A06C26110003C0A05018040004018100809000080A050281004030380C0",
            INIT_RAM_3A => X"5A1C75AA9F2C8BBB5AEE1793D9AC9B41A0D088C46231188B46231168B451E0E06E339651",
            INIT_RAM_3B => X"E6D3D299B2F66C3D9749D5837228AB37B31FCCF9AA5592DB54A38FA6C140180E0A058342",
            INIT_RAM_3C => X"6050281406040305C2A0F0B0382C0D0602C04020201C0A2A1A9147C441A0CC562B178480",
            INIT_RAM_3D => X"A9449A08F06F339207C2F0480802141307428110483C1E050080804010301006030180C0",
            INIT_RAM_3E => X"6580300012040A85C45A2CBDEEA12C87B919CDF73B718EA4462352A954EA553A9D4EA752",
            INIT_RAM_3F => X"C441A0D47624188680AB24829D2ED560BA0D9318E26962BC7FB9DB4F072AFDCCBA48A243"
        )
        port map (
            DO => promx9_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_9,
            RESET => reset,
            AD => promx9_inst_4_AD_i
        );

    promx9_inst_5: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"6030200400060201408040180804020283C3C08040781E0E088100402030243E1A1B920B",
            INIT_RAM_01 => X"A9D4EA753A954A251288B45204E068338540A020D07808101387848020602C1C00048000",
            INIT_RAM_02 => X"2E277B653C3B15244A061008780A1A0309C47A2CFDF2A1348BB9196C260AC56C9C462352",
            INIT_RAM_03 => X"40400034402B1F940AE451AADC9834198982EBE6241DB4F066B19590CC53BE90B155C158",
            INIT_RAM_04 => X"C1F0080C2E250A02C2611078140401030180A05020100A050783C22170805C2E0E028100",
            INIT_RAM_05 => X"EA653A99388B4223528954A251188B41A09047A3C9C0DE762A88C3835260EC6A00100582",
            INIT_RAM_06 => X"B35A3BA9935882C41C0EF67B3612924E9F10A4F018542C2C0F06407A2CC612B33D8FBA97",
            INIT_RAM_07 => X"82513014060707030040507830302D24180A0482895C80551E0BC344F675DE42E56DACEB",
            INIT_RAM_08 => X"A3E271147A35158F0742C1D8E87231140983813090400802000180E06028100605030049",
            INIT_RAM_09 => X"7A2CFDF2B1358FB9D488D46A51188B4222D068341A0904813C9E4E2703798106692B9387",
            INIT_RAM_0A => X"005603E9FD2D7E5C6D34451C7641077ECD246C57630A3CB4599C0B417018144E36110E05",
            INIT_RAM_0B => X"C06030180A021113C6212219288A260201C040300034263B391E1566C32028C0580D0B40",
            INIT_RAM_0C => X"06F2C9BD0C622495C925128130602F239188C462291078421D0C44E2D0A0281C0C0101C0",
            INIT_RAM_0D => X"20B0A8785612239A487A2CC5EEB13C8E351168441A11168341A08F6823C9C4E271381A0D",
            INIT_RAM_0E => X"A853E8B4E2053C81C16066BB9DB10AC043A7B2B9AE1A8D5F6AD1DD91B6AB495E94449B43",
            INIT_RAM_0F => X"0161286C120D018000C070301C0A1E200CC964B248C8802E1380C02010002C14372C1BD3",
            INIT_RAM_10 => X"271381A0D068341BCCE652EAC902732596CB65B2C12000392893C90482401C7A3D220C44",
            INIT_RAM_11 => X"F026638D10A832954000D028448C57229A555A2CFE12B133852E8E67A3DA0D088B411E8F",
            INIT_RAM_12 => X"8040300C0025242A982D2919710A760001C1C0106B81E719964AE451E7C436771B973CE9",
            INIT_RAM_13 => X"44E2293C7C331989C32200F0702016018000A0703800024D2488C9642208AC74311A8840",
            INIT_RAM_14 => X"47239A0D047A3C9A4E068341BCCE6733178BA552B3596C5508934CA6D3386808542A9889",
            INIT_RAM_15 => X"D0A9E249BD165B2AD1AA85AB84FE662F8180414030B0AC6047A10D399C863AD3387A248F",
            INIT_RAM_16 => X"84B1C8A4563A188FC460C0280C102D2524642D6942993C2138184DD7117A11B5198D5F9F",
            INIT_RAM_17 => X"22E1E008507F3D158DA5C2D1247E421886442180E8281E06060000C07000144E7512050A",
            INIT_RAM_18 => X"189C863EE33A611C4E2723D1E8F4783419CCE5F2F178BC562A954A84D24B39884C0C0B82",
            INIT_RAM_19 => X"69B5B16914DE75C660A9A39194926023140CE66528B8A6450400C0A05138F4D85D3C1401",
            INIT_RAM_1A => X"E070310C2E6F339B8DA4C2190864331D0C45E1A0683C2804201E220CA6725CC61B411F8B",
            INIT_RAM_1B => X"84B229BD9C8F291E8B4BD61E99B6A248A010E7E3513C7C3B198A8401F0E044000E018180",
            INIT_RAM_1C => X"E131187876AF42812AF88C463EFB25489C4D271389C4E06833978BC562B158AA55269349",
            INIT_RAM_1D => X"95087AA0FA672F1407C45049B4A0053896CDE572A91CA62D2981072291D04C8E14018100",
            INIT_RAM_1E => X"42F0C8200C04008180E07518546C65301D8CA60158EC78431D8E8723116830020E238F8E",
            INIT_RAM_1F => X"C552A9549A4C2212C864323105DED54EA857ABB753D998AE5DA65228D39978782F1008C8",
            INIT_RAM_20 => X"038128340806020080C03048908475392CA7F80C4632CCE1389A4D269389C0D0672F178B",
            INIT_RAM_21 => X"844228081004021B17AF1AFABD469365149BC4F2D0C8040301070683C218EC76280D9088",
            INIT_RAM_22 => X"ABB8F1E4A83C1A0F08225098200C04038040E06270EC44422A114AA4D269348A4D271349",
            INIT_RAM_23 => X"269341BCCE5E2F158AA552A934984C2590C86431D0CCF2DC7CB49E4F274385D70460BE93",
            INIT_RAM_24 => X"80D030382A15120742203020100A04020180606038204623191EDD188C860680AA38180D",
            INIT_RAM_25 => X"845239389C402B1388C451E0D0180400929E0DFE355CE084308446A131A80802040200C0",
            INIT_RAM_26 => X"6FD96426D2F279AA9FCBD58238D0462508C6E240883C0A04008040E0542A1440320F08C7",
            INIT_RAM_27 => X"189CBE1A588138180D2683799CBC5E2B154AA552A93096442190C743A1C8A094E173CD61",
            INIT_RAM_28 => X"616018040805028140A030200C0607020100A04028180E07028100604030382229158E4D",
            INIT_RAM_29 => X"2051119464130306C0E451C00CC0492D164A2502B9388C260E1B167BA7F9D8D449029101",
            INIT_RAM_2A => X"432188B46CCC78B69BB279FD2AFB3E61AD584A14BA249053140A05A1A0483C0A03020840",
            INIT_RAM_2B => X"40506058101A020003391CFDEE26703317CC0603399CBC562A9549A4C2611086431D0E87",
            INIT_RAM_2C => X"AB89584000050601C1C040181804020F8845E27128583A1A020080A0502010000F020100",
            INIT_RAM_2D => X"6020801C0A030200C0801013248025000040C140698CC86A25174E6622E9B8020700935A",
            INIT_RAM_2E => X"A4C2590C863A1D0E46229148AC4293813BA47779B4A713618338A3C82341747843160C03",
            INIT_RAM_2F => X"4160281800080301C0C02010140C111086845A2D35E1F47733158BE5F2F978AC552A9549",
            INIT_RAM_30 => X"E8646A08CC510D00882A53C358F660060140A060300046210207048071A8702A240D8602",
            INIT_RAM_31 => X"2953B22878341D0DC5C1A0481C0A0D0600C0609001080454318086A7D3D8F4D45312994D",
            INIT_RAM_32 => X"A552B154AA552A130984321908743A1D0C462291408842347542EE15F9A37A5507703A91",
            INIT_RAM_33 => X"814020744C1312090381B138140C01048140606008100A070B05079ACD7E01E4762E958A",
            INIT_RAM_34 => X"E7534210D08040205086B58AB50259150180E06010140C05030080E030084C0A010F8044",
            INIT_RAM_35 => X"F12B7D027B259541DA27F3F998CC4A3808450240383804030601406001810026230DA3C6",
            INIT_RAM_36 => X"9B4D8601F6772F154AA5426134AA552A130884321908743A188A452281009C3A1C22AF65",
            INIT_RAM_37 => X"C181A01C2C010B83C221F048542C0B0A8744A1A090402001000001E060280004040601C1",
            INIT_RAM_38 => X"A100219C78223F004A08149268BAAC51890924565AE54877188180C07030180A040301C0",
            INIT_RAM_39 => X"0201387C34170E0E13D31AD54E2F338AC81E6C43B134AE4C1B1108813020280001030340",
            INIT_RAM_3A => X"0000300C0E060100C09ACD8E2A047033178AC562A130984C2590C86431D8EC7431148A45",
            INIT_RAM_3B => X"E06038180E07038080E22058900C000804832100701400090986C3A1D1105C0411048140",
            INIT_RAM_3C => X"8040100000030281008040481C6C581815D12955A29E5A7E692F99EDF512AD6A8B1C0180",
            INIT_RAM_3D => X"63B1D0C86431148A040270F05C3E1304898A87376CF2491877BA5F8CD3D9C0A05F2499C4",
            INIT_RAM_3E => X"4140E0683411000040402038180C050301C07ACD4632367832954AA4D26130884C219108",
            INIT_RAM_3F => X"CC76B3254477310180E070301800070381C7C1808850021006804201603054000A080302"
        )
        port map (
            DO => promx9_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_11,
            RESET => reset,
            AD => promx9_inst_5_AD_i
        );

    promx9_inst_6: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"4BB3819CC4582F0BC360B0180C040306850180403800D06D149A53CBC5437656F65D5D98",
            INIT_RAM_01 => X"84526930863B1D8EC763A190C45228100803E170B0582C0F098244A3C14911E512833B25",
            INIT_RAM_02 => X"E0F0881006100102C240C0E07044100180402010001C000201818079ACCE267C903210C8",
            INIT_RAM_03 => X"1046ACD26F5F6F36D470C40A9D3687080140C000301C080503850860903000200F0C0402",
            INIT_RAM_04 => X"21B0C82836133432194DA42170CA67158A02A1D020301803018182C0E050148E5E5C39D3",
            INIT_RAM_05 => X"592C9652C6C13610876442210C7432198EC7432188A4522F10064341B0A04C1602018181",
            INIT_RAM_06 => X"80F090580626030181C140400808020585C141D0B0944C3B110080207000080604008482",
            INIT_RAM_07 => X"E0A0081472603A4D58ABE9D425FD3070561D0EB7A2DD3228000100A06028140E0602A046",
            INIT_RAM_08 => X"0111006430170404428260D00C3C140902C062B1107C06002A10C6A27040740C070682C0",
            INIT_RAM_09 => X"A02028100A00060082392CD67AF9123A92C86431D8E86432190C86431148A452220E05C3",
            INIT_RAM_0A => X"E07020140E06029EC36020F0D4601C08828140401014260A0283808250E8984C290A8080",
            INIT_RAM_0B => X"C2A0B03C1A00090241E0F0501C3EA63CA5936BF9F35DA2FA7A43DCB1175AC0C60A0B8500",
            INIT_RAM_0C => X"431148AC3C080D06C462B150A4321A09068361F1786C2E2F13854260A0481C0C09320E87",
            INIT_RAM_0D => X"6130A89C6E251103C160503828000C048141389C9667154D4796C8432190C8622A190C86",
            INIT_RAM_0E => X"2F56CAB81A1B050441006030140001018E424220F0DC720F0D91130050B00C0C111784C2",
            INIT_RAM_0F => X"80B0B00012322E0C04C290F0281A1F0602C0E0105030262C3B9F528C487F3220EA7D3E1D",
            INIT_RAM_10 => X"432190C86432190C86429128843624120705A2C1188C461A0E04C3C28148A04020138582",
            INIT_RAM_11 => X"2030800022040700C36160F8BC5037160100C03068544817000184188C564B2D6C609CC8",
            INIT_RAM_12 => X"0E2774BE58AB8BC65EAD8540902A0B058241E07000380A05018F470120F80C341F058D01",
            INIT_RAM_13 => X"028150A85A18100981A120A80402702B12C74250E07446140F0744A1C0A8343C2825A511",
            INIT_RAM_14 => X"389C4E4B31889A2109432190C8663A190C8522C158B85A25128944A2C0E0504824120984",
            INIT_RAM_15 => X"838290904C010F0542A11000140E050E0282207140A452281A00C10190F83802150404C6",
            INIT_RAM_16 => X"C1F100BC50301C0D44C9A56AC1C6F97B361CE8C0900818140602804080482410060B8B06",
            INIT_RAM_17 => X"A1D0A0503A1D168984429150A86C1D0F85C4A0301800127B31174741D0F8A05815100DC4",
            INIT_RAM_18 => X"0241F8F86A36028F4859AC964F459CAE324E642198CC763A190C4542B100C06E37138984",
            INIT_RAM_19 => X"40B0D848120C128980C141F03054190A00444311F8F4081610800341E100A45431178640",
            INIT_RAM_1A => X"830108D84A1B218F0AA53250EC843A208F8540164C324F2F780711C49130984E0F028502",
            INIT_RAM_1B => X"039198C86231148C05E270F0985820178846431118AC54281009C2801008242E733095C7",
            INIT_RAM_1C => X"A25100A8562C158901A212812CC658228B467A3CD66F479FC2C7D3E5B218EC763A190A45",
            INIT_RAM_1D => X"E591A86C2A070382404120584814130D84438400D06098290D084421D068681415068202",
            INIT_RAM_1E => X"C1A0884008514A1A4924C210EC923C27964F06B2A958DA64291184A0F0001C320D2797C5",
            INIT_RAM_1F => X"885298E86432188B05E341E0EC742A150A4522F100AC6633180A4462C160D06422138604",
            INIT_RAM_20 => X"A350384808101003C02050C8AC5A35168C01C240D990C65B2D98CB9A3D1E8F479ACA585E",
            INIT_RAM_21 => X"40C068100C042A9344647058601E050F000181C0705016032F0DC721D0289062090D8AC5",
            INIT_RAM_22 => X"A2E198B46A2D150A048090503C16A248A0CB8632D168C25F299D11AA2422810C6D328B86",
            INIT_RAM_23 => X"5A3D1E9347A3D062EA0EC3E9086432190B47E501F8F46833150A852210A8D878351D0B07",
            INIT_RAM_24 => X"82B0D87048200E904264200094340C480806E22140705A361A8B0424633A3D0C6F3C210D",
            INIT_RAM_25 => X"2D6572CD3E732912C441C018080605250F4A60E0206836130482C2614098503414129187",
            INIT_RAM_26 => X"42314940903A170305E47239187E3D198A85C230802002126F2FD628F439F8EC764429D5",
            INIT_RAM_27 => X"480389E0E6893CA25139ACD66F47A3CD67EF345691D0863B1C100C6622811C6E361A8D05",
            INIT_RAM_28 => X"40B07090301B0708C8A2F0B0C410490C88C640C0A13C76C20283464050E0D45A36208402",
            INIT_RAM_29 => X"ABC56AB176BE7FBCA311372AA50C6B2B0B86E0C01008020B299144C22028043C090A0682",
            INIT_RAM_2A => X"E7C2D12070381F8D876351E96CCC3A1D818524929160A04E1A0844C2A048282C5A7BCBDA",
            INIT_RAM_2B => X"433000006869270C0205835A111A94401750399CCE6B259ACD6672F7F98AC0BA441F1791",
            INIT_RAM_2C => X"C2908018101504848240B060303611000B8503A38098724A0D8B45058080646E61068480",
            INIT_RAM_2D => X"E1B090344A7652456391569492531887C063ED06616CB85A278EC420202008023A1F8B03",
            INIT_RAM_2E => X"38CB2B789A44229E9428E3616CA442208DC7836239B4CC4226028964C2A16CA24F1E88C5",
            INIT_RAM_2F => X"4190A9044A172387450884D904A45D378D8948B412151A9C681603399CD667359BCD66B3",
            INIT_RAM_30 => X"E0606008025A1B08C0C07000082C1F01058380B0E8703815149149D2E2498488501F9ECF",
            INIT_RAM_31 => X"C6633170A441278D4442506860746F5325A5107E76D6993C9FC60C6B43A0F0B85E198AC1",
            INIT_RAM_32 => X"599CD66B359ACD66B3594B2358AA4C1C25564973A954BA5D299408A43309FCBC3F298A88",
            INIT_RAM_33 => X"E4D108B84817108EC98031681C3E161F9486C1249128D66331120004842299489F56BBEE",
            INIT_RAM_34 => X"E422609022551E8040806020000A4E0F89428110482022110B80016140F0744C2312A885",
            INIT_RAM_35 => X"6783D1C0B27F24140E26934198B84A208DC5828110F8664858AA5571E78489DCF8B78810",
            INIT_RAM_36 => X"61A3F3320ED5CCBF1E39ACCE673391C8E6B2F789E23CA83B18255769244A25027A512BD2",
            INIT_RAM_37 => X"612068943A2512940DC850EA9037463D0D01A2B3C96C8EA80C878424D251B9149A2A9C41",
            INIT_RAM_38 => X"AE989371DAA7190AC8213050581C04020100E050200C625A190F848120606C382A078243",
            INIT_RAM_39 => X"0D281C8A23018540206B94B904C680351CCF67A391A4CC4D1D8A05C2B0F8B8060145AC94",
            INIT_RAM_3A => X"44C2F1ED5E873B818000007A71FCB1734E1D399CCE472599C8E43175C6E930863B1A2199",
            INIT_RAM_3B => X"4130E050460310008201107814380C088747046549005E553311038732C8507A2D130907",
            INIT_RAM_3C => X"02D1481C18041E30196973A9509A442389C46150D0000E05028200E0503008DA491A8503",
            INIT_RAM_3D => X"B283693076341D96159079C57EA72A883E1C0ED60A0CF67442A351C9E4A1C8D4672B10C7",
            INIT_RAM_3E => X"230009B0561C0909C8A642F9ED307E3B8641C0B000054EE78FC629399C8647239ACCE7F1",
            INIT_RAM_3F => X"A0602814B234208DC1E040380436010482C2E05098400C2008811484C21098C4423719C1"
        )
        port map (
            DO => promx9_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_13,
            RESET => reset,
            AD => promx9_inst_6_AD_i
        );

    promx9_inst_7: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"E9853A39086B30158A44110808100E03A05BCC560B38F2270F04C2E0B0602C160A088040",
            INIT_RAM_01 => X"391C8E472391CD69F030422910763D23908F51AB15C6C92B89C2A07087B1E8CA843FA414",
            INIT_RAM_02 => X"4212F8B4C4490F2305ADB0E914905421104AC683F2A900710C0782403018000E86593D5F",
            INIT_RAM_03 => X"40A0982C1614090000E01020047C151E8580803058305E0A0A88C22041103C0A100184C3",
            INIT_RAM_04 => X"0DA821B09C817226988E35E36DBE96461C0B44405028220F028099706540DC40270A8701",
            INIT_RAM_05 => X"A1D01810000254AF94391CCE47239ACD68310FD26930763C2310090B19558AD15592449D",
            INIT_RAM_06 => X"E040385C30070283C46E72A96D2A4523114CE420A8B8926A53860AABD59A395E841D8C03",
            INIT_RAM_07 => X"003160B45C2D170283C06008402A020C00802020485006361E114663A0108830030B8102",
            INIT_RAM_08 => X"24D4ABDE91468E45570A248AEDA6D27BCF30552B6BD604C157A48E4350982C2409070182",
            INIT_RAM_09 => X"2D05FAF5762D220E85E2205010060002319459ACCE67339ACD6631D2832930883C229188",
            INIT_RAM_0A => X"005090845808188800E010201C1C01000141E1448AB616961F9AC3667291A4AA6E3A3197",
            INIT_RAM_0B => X"A1F1283034090401870010D88076240D05816000404C06070001C08130605C0C3A2E8D04",
            INIT_RAM_0C => X"55F57974863B1E0F48C40279C566B152A04DA62252357AB75CB8590C26C335F8EC6D2ACB",
            INIT_RAM_0D => X"A555638D38BE59B85B6EF5BA304256271108234128500A0E00050059AD1667339ACD6671",
            INIT_RAM_0E => X"00B028502C663913402050C8D4100F01048442513874302A2280C762A03D110AAE2F1F87",
            INIT_RAM_0F => X"486349548C3B210B84E20178743812078086805168C4380004040101202058120A0381C0",
            INIT_RAM_10 => X"59ACD66B4599C8E431B698499CBA441D8F07A461F900804125148A450279187A31272754",
            INIT_RAM_11 => X"0031500AAE4276539CCF542B5572EE93309C08B34960C46623130943E138300A06078201",
            INIT_RAM_12 => X"C0E0881C1810050402A1D0B86C006E331369007068681C080F05C421B05850122B1A0D01",
            INIT_RAM_13 => X"C46228F06834199D54A903595C8C45218E8683A1C0BC3A1B069A43A220F8483C110303C2",
            INIT_RAM_14 => X"65D1A8340C0F078002599CD66B359ACCE431D70A7395026E26110763D1F1188E47201008",
            INIT_RAM_15 => X"2290206C52260F03C180C1580810A09F3DDB90273B361EC86833DBA84429ECD4612D1DCD",
            INIT_RAM_16 => X"227020184A0F0A82C10030683C320209850240C0D8604EAA009945A0E2503C34280C8885",
            INIT_RAM_17 => X"C4D220F478351E0F47A341E0EC6633199013CAB461BC8A441A0F49C56321044E1D0E8C84",
            INIT_RAM_18 => X"C8C0E9D90094399E50866220181C08088442398C8E47239ACD6672186B8D2A0AC1521E4C",
            INIT_RAM_19 => X"C35218501009158CC522E1A864483826854482E1B80C0206168D068813A885E8BA569FD3",
            INIT_RAM_1A => X"C52391E0C234251104A1006838420209848060C098240E110D05C261F148DC36B31796CB",
            INIT_RAM_1B => X"390C35F2C75BA84C96265220F0783C1E0F07834198C856331A0B4DEB6541ECB04521994B",
            INIT_RAM_1C => X"ED649B3194C05B25CD05F2827D2E8E4E25CE463168140C0F040442188C4647239ACDE6B3",
            INIT_RAM_1D => X"8220180C280541A2C5C3D040AC66290C8AC622E2B1545410020C8003E1F848040025144A",
            INIT_RAM_1E => X"0AF55254D45921158A05E4FAB52A40361B476110203C1A06038340E12030582C3F000202",
            INIT_RAM_1F => X"D7FC3E031191CD66B47A2C863F0F7FC2DA6005D218EC783C1A0D07633198AC562B158ACA",
            INIT_RAM_20 => X"2471E0282C1F2AA21524337A8D90914F0ACD468059F92EA058A082834128340C08080442",
            INIT_RAM_21 => X"60D04008162B0E008362D068D00C075A19D2E67190B88A37230B454251B0609049A51646",
            INIT_RAM_22 => X"633198CC5633150AC667F602E8D6883B16CB4764FA8CFE551A9B89604109B0228E118740",
            INIT_RAM_23 => X"00C020181E110C044396DBB5FF0F8FC4E4B37A2CCE431F87C35F24065220EC683B198CC6",
            INIT_RAM_24 => X"E361C981D4AA30B44A2301C0181A034937150861630D9F405400526043B2312AA24B9E83",
            INIT_RAM_25 => X"24B1408402DF138314A15080BC3A10040304A25018B8041A020A4F27F1B92086542209C5",
            INIT_RAM_26 => X"E5D1D8EC663B198CC6633198CC6633190CC6A394F3553CA2471A4AE5C3F2510E53260BC9",
            INIT_RAM_27 => X"EE908960B89E39800700C0303C1010088643553B25B6FD7FC3E27259BD16672188C7E124",
            INIT_RAM_28 => X"E271B0CC9E310E09C66197FA70F87933A54D64A210EC1E787AE61EB915395918C897FFBE",
            INIT_RAM_29 => X"075311AD0C5C699AC9A4F3D9A03E350988126C50685C38390B8E014161D8A824081FA20D",
            INIT_RAM_2A => X"392CDE8B3591C86124C54218EC7633198CC6633198CC6633190AC542A2A2A5CEBF58A3CD",
            INIT_RAM_2B => X"319C26C190FD7611D38853799CCE6A2B04418050283C2C090C868434AA9592C96DBB5C31",
            INIT_RAM_2C => X"E0D298F86C2F2609D5E6D32940C26B1B15D565C342412CC048B9CE654299342415712A54",
            INIT_RAM_2D => X"62B1599982E166B19989C57A1942863D9ACE053221309AA44A24086DD131B0867B179008",
            INIT_RAM_2E => X"141A956AB55BB25BAFF81C966B359ACC6365E54218EC663C1D8CC6633198CC6633198C85",
            INIT_RAM_2F => X"A662F1DE564A51C7678E7512856A72BC5C954A746224F24F020300A060783C22190C8484",
            INIT_RAM_30 => X"4A2599BC82661C0D4FE902CA9D6E9D3D18580B73AB49E64716A8422963CA35808C58244F",
            INIT_RAM_31 => X"633198CC6633198CC6633198A8A8B970329A2CE5F22120A093B78EC7A1D158A431219ECA",
            INIT_RAM_32 => X"C070805C20190C8683149A554AB75BB1D92DB77BC6031189C461E7E5C220F0763C198D06",
            INIT_RAM_33 => X"08459AB97CBB56AC0E0773542D2F798F3EE60B1BCC4AF60C7C2494C9447988A8270E0341",
            INIT_RAM_34 => X"6892914CB63524A89A29631988BE412A9B07680441548CD24D9F106C142208E6543B1540",
            INIT_RAM_35 => X"26C220F0783C1E0EC6633198CC6633198CC6633198CC5C3D533D616E75C2E19513692152",
            INIT_RAM_36 => X"88B4494C5A06028381E1008860221A0C86C4148A554EB763B1D8EC96EBBE030F87C3DE28",
            INIT_RAM_37 => X"D0D2620550070094C26A3AFA09E0E071A8D368B498BCA251AC3E4E52E752AF0DBA2E9FD2",
            INIT_RAM_38 => X"B268DBE5B0CA89B95CAA2439D8DC7C2F388E879030F90C792B264E45E4D0D0E8B257A790",
            INIT_RAM_39 => X"965B75FF0180C3E02747D22110863B1D8F07633198CC6633198CC6632158CC562B169BDA",
            INIT_RAM_3A => X"76EE23E926AA542448C6E1E0200C0E0785C101808868421B120B05149A8D2AA55AAD56AB",
            INIT_RAM_3B => X"A704A2E952B6A0ABD2C836C2615E47268E8C8EC88C3A63006F4B546841A8E41B42643E69",
            INIT_RAM_3C => X"633198CC5632198D878AE8BD4AED338944DDABC40A1CD4F140230B2CA121D83C6C2889D2",
            INIT_RAM_3D => X"551A8D269552A954AA55CB35DF0F80C3E0AACA522110763C1E0F07833198CC6633198D06",
            INIT_RAM_3E => X"8372693CB64C995C2ACA15723156823F1A4720D0281C1E0F0B840221A1108C4624160B05",
            INIT_RAM_3F => X"EC46B398EA71299DC8E845730D56A359B79C66301CD98D8F7BDF140B2B248A79B174B515"
        )
        port map (
            DO => promx9_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_15,
            RESET => reset,
            AD => promx9_inst_7_AD_i
        );

    promx9_inst_8: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"1C0E080492490092512090492512C964A2592C92482391C9048239208E4A24924944B259",
            INIT_RAM_01 => X"1408040281C944A2491C8A0402820924923114080503124944A2411808050281C1009238",
            INIT_RAM_02 => X"6E371A8BB51A491482411C8E4724124D14823D188B451351A8D46228924724124944A239",
            INIT_RAM_03 => X"24924A26928984C25965B5196CC65B3198CC66351A8DC6A30D66CC6A33188B361B51B8DC",
            INIT_RAM_04 => X"20100803820124A249289248251249049249249249241208E472391C904723920904A251",
            INIT_RAM_05 => X"2C904623120944A2391408040281C924A2491C88030281C90482301408050301C9048241",
            INIT_RAM_06 => X"6233186B359B31A8D46A371B8CC55A4D14823D1C8D46A351C9047A391A8B4512C9A8D462",
            INIT_RAM_07 => X"180E4824124904725130964A261289A545E759AED88D46E33186BB6233198CC662ED66BB",
            INIT_RAM_08 => X"180C070412494492592492492411C924B249249248241208E47241208E47239180E47239",
            INIT_RAM_09 => X"3514492412C988D461248E4502920964B23914080502818924A241180804028180C47030",
            INIT_RAM_0A => X"5DAED88CC622ED66B361B0D76AB55AED98C461B3198C455A6D2482391A8C45A351C8F47A",
            INIT_RAM_0B => X"188C47239209047241248E4724124924924924944B28A5524B4DAE5DAED98D46E33176B3",
            INIT_RAM_0C => X"180C060381C0E0824020904825128964B2592490482411C90482391C8C472391C8E47239",
            INIT_RAM_0D => X"451C8D462311C9048A351447239309C8F461288E4502820964A23914080502818104A241",
            INIT_RAM_0E => X"5DB0D98D46E33166B355ACD88CC622ED66B361AED669B51AAD56AB55AED98BB55A8D369B",
            INIT_RAM_0F => X"100A06031180C4623920904723118104823924924724124964825934AE996D34965B9DEF",
            INIT_RAM_10 => X"100A060391C104A2411C0E0703820924A2492892492492492482411C8E46231188C46028",
            INIT_RAM_11 => X"55AED88C45DAAD46A34DA08C4622C9E914923D1447241311E8F461248E462301C9449231",
            INIT_RAM_12 => X"65B6DD6D3CF6DBEFF75DB0D98DC6E33166AB51AAD76C461AED76B35DACD569B49A8D46A3",
            INIT_RAM_13 => X"1C8E47231188C06231188E46039188C050311C8E472411C8E47239180E482492CA4984B2",
            INIT_RAM_14 => X"208E460281812492411C0C070402090492412492472392092492411C8E47239188C46230",
            INIT_RAM_15 => X"55AAD46934DA4D46A355ACD98DC6A2ED56934DA28F451289C9249B411647241351E8F459",
            INIT_RAM_16 => X"208E4A27A65B4D74E379C0EBBAEDF7BFFFF75DAED98DC6E33166A351AAD66BB59ACD56AB",
            INIT_RAM_17 => X"180C47230188C06228140C462301C8E47239208C050311C8E46039188C060311C9047239",
            INIT_RAM_18 => X"4512452392C9A8D2592490460381812492411C92492412092482412090472391C8C46231",
            INIT_RAM_19 => X"49A6D46B35DAAD469B4DA6D268249A6D56AB55AAD98DC7230D368A4DA8D2462249A926A3",
            INIT_RAM_1A => X"180A05030140C0724138AE986CB61AA954E381EDB2DBEFBFDFEFFF5DB0D98D46A331669B",
            INIT_RAM_1B => X"188E47231188C46230140C06231188A06028140A06028140C06028140C05031140A06030",
            INIT_RAM_1C => X"51AAD466A209691492411848251309A4F2612894492492494492412090482411C8E47231",
            INIT_RAM_1D => X"5DAED86C46630D669B49A4D46B359AAD368A45229148A4DAED96CB59AAD98E47230D368A",
            INIT_RAM_1E => X"140C07239188C46231180E460281C14514D36132D54AA6134D84CBF7EFB8DFFFBFFFFFFF",
            INIT_RAM_1F => X"1C8E46231188A45229140A052311C8C46239188A06031140A45020100A05028180A05028",
            INIT_RAM_20 => X"5DAAD76D46A2ED368A51ACD5482389A524A2491E8D27139208F471309449241209049241",
            INIT_RAM_21 => X"DB75FFFF7FFFFFFFFF59ACD76C361AED56933D20936B35DACD368249A6D048255B51D8DC",
            INIT_RAM_22 => X"209047039209047028140A05031140C060311C8E4D2AA5530D84BA592C9A6DB65AE965B6",
            INIT_RAM_23 => X"2C90482391C8E46239188C46229148A45028140A05028180C46039188A050301C0C07249",
            INIT_RAM_24 => X"4DA6D368A55B51D8EC61AAD76DB7636D96BB61B2D96AA4D26954AB55249148A41208F46A",
            INIT_RAM_25 => X"6132DB6B269A6B3DBEF7FFFFFFFFFFFFFFFF51AAD66BB5DAED6693391E946BB662ED368B",
            INIT_RAM_26 => X"1C8E4924928944C2713C984B2592C984A261349648230140A07059412C954C3592A954D3",
            INIT_RAM_27 => X"51A4914823D1C8C251208E46231188A45031188A05031148A05028140A45030140A05028",
            INIT_RAM_28 => X"4522D46C36A331669351AAD468A51B71D8F46DB2DB6FC86431F8EC763B1C8D361ACD76B3",
            INIT_RAM_29 => X"592C954AA5D30D86B25D32D84BA9E65B8DF7FBFFFFFFFFFFDFFFE74DAAD76C46A35198AB",
            INIT_RAM_2A => X"140A06230140A07039249A5752CAEE7B3D8EC767B2D96CB53248E3489C4D25930A4974BA",
            INIT_RAM_2B => X"76391B8CC5DAAD469B49208E46A3096492391C8C46228140A04020100A05028140A05020",
            INIT_RAM_2C => X"4DAED98D46A371B8C355A4D46C36632D76A355AED76B35DB8DF90C7E41219148AC5608F4",
            INIT_RAM_2D => X"BEE36CB0B2C984F28A512C964BA592E934AA5D2C997CED773BFFFFFFFFFFFF7FBFDF8DD7",
            INIT_RAM_2E => X"140A05028140805028100A05030180E492D2BEE5B2D8ECF63B0B8EC2DF71D96C765B1D85",
            INIT_RAM_2F => X"92C561B0D86BF1C8D4622ED56A349A29046A31164B251249047239188A05028100A04020",
            INIT_RAM_30 => X"FFFDFFFFFEB75DD6E355B31B8DC6E391D8DC5DA6D36B369B4DA6CB61B4DB6DB72412191D",
            INIT_RAM_31 => X"BAD96CB6DB6DD6EB7DBEDD6FB86BED9594812CA0564A24D28924AA5528BBFB6E7FFFFFFF",
            INIT_RAM_32 => X"188C45031188C05028140C06028140A050281408050281C28B3D96C75D6EB75B6DD6DB65",
            INIT_RAM_33 => X"7A3F20904824322B1D8AC3608EC6E33176B351A48F472391C8B259289249249208E46231",
            INIT_RAM_34 => X"2CEBB7DE7FFFFFEFFFFFFDFAFBEAABEDD6E359B51C8E46A3B1D8E469AED66C36DBB1D8F4",
            INIT_RAM_35 => X"BAD96DB5DAED76CB65AED76BB6DC2E16FB6DAED96CB75C2E36FB8E92244F2814D229249A",
            INIT_RAM_36 => X"249048239188C46231140A05028140A05028140A05028140A05028140A060398E63B0B7D",
            INIT_RAM_37 => X"72391B8E47E412190C8643219047EBF1E8F4763B1B8D461ACD469B49A08D4622D168B251",
            INIT_RAM_38 => X"C2D75A440409E534A2CF6FBEFFFFFFDFFFFFF7F3BAED375B0986CB61B71D8F4723D1F8F4",
            INIT_RAM_39 => X"140A0836DCB5F6EB5DB2D76CB5DB2DB6BB6DAAD76BB55AAD56AB5DAAD96AB55AAD76DB75",
            INIT_RAM_3A => X"451E8D45A2D164B249209047231188A05028140A05028140A05028140A04028180A05028",
            INIT_RAM_3B => X"6E3F2191486432291482411F8FC824320B0C82C15F8F47235198CC6A35198C459AAD369B",
            INIT_RAM_3C => X"AED56AB4DA65128944AACD1B6A234986EBA6E37FFFFFFFFFDFEFD6F7AC9A6BA552A964B2",
            INIT_RAM_3D => X"100A05028140C060301C906FB8EBAD96AB55AAD76CB65B2D96BB5DAED76AB55AAD56BB55",
            INIT_RAM_3E => X"59AED76C359AAD3693411C8C4592892492411C8C46231188A05020100A04028140805028",
            INIT_RAM_3F => X"30AC944AA5526964AA824764B2592C963B1D86C160AFD7A3F1E8F476391C8D4662ED66AB"
        )
        port map (
            DO => promx9_inst_8_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => promx9_inst_8_AD_i
        );

    promx9_inst_9: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"C2D76FB85B2D56BB55AAD569B4D9E4D248EB511E5029244EBB6DE7FFFFFEFFFFBF5B4D2C",
            INIT_RAM_01 => X"100805028140E050301C0E4824920904925128ACB2D6DAED56AB55B6D96EB75B2D96CB55",
            INIT_RAM_02 => X"6631188CC5DAAD56A351AAD66B355A8D167A39188B241208E47231188A45028140A05020",
            INIT_RAM_03 => X"FFFDFEFEFDB6BA893C75A24E28938985449A8EC965B258EC763B1586C15E8F472371A8D4",
            INIT_RAM_04 => X"AED56AB55AAD56AB4DA6D369B55AAD56AB55A6D36793C8A38D347134984E2A2C2EBBFFF7",
            INIT_RAM_05 => X"140A05028140A06030140E0704120104925930A05129A44A2524AA6DDF6DB5DA6D36AB55",
            INIT_RAM_06 => X"7A3B1C8DC6A31176B355AAD56B355A6D36934926D56B359A4CF46A2C9047239188C46231",
            INIT_RAM_07 => X"349C6ABA6DB7DFFFFFFFFFF8DB6BEE16FB8EC76371B96D338D548992C562B0D82BF5F8F4",
            INIT_RAM_08 => X"BEDF6DB5DA6D56AB55AAD76BB55AAD369B4DAAD569B4DA2D168B449E4B218D3451C4D271",
            INIT_RAM_09 => X"208C46231188C45028140A05031140C0603920984F2925938E2944B2DF6DB6DBADF6CB5D",
            INIT_RAM_0A => X"82BF1E8EC6E351B8DC6A351A8CC622ED56A34DA2D149345208E4723D1E9149B49A28E451",
            INIT_RAM_0B => X"7DB0D1471389C5028944E9B4DE7FFFFFFFFFEFE9ACB5DAED56CB5DB2DB6CB75B2E16FB75",
            INIT_RAM_0C => X"CF6BB7DBFD75F6CB65B6DF73D75B6D96BB55AAD569B4DA6D369B4DA2512893C9A4D2591C",
            INIT_RAM_0D => X"24964D47A3D1A8B2491C8A46228140A05028100A050302018512B275C72AB75BEDD6FB85",
            INIT_RAM_0E => X"AED96CB65B2DB6EB8576391B8CC6233198CC6230D66B355A8D368A3D1C8C46A35188A251",
            INIT_RAM_0F => X"9E4F2793492471D6BA451E502894924954AACF6DBDFFFFBFFFEFAEC2D76AB44A2536AB5D",
            INIT_RAM_10 => X"C6E1B3DAEDFEFF7FAECF63AFD6DB2D368944A2576DB7EBAE1ADB55AAD56AB4DA6D168944",
            INIT_RAM_11 => X"3114492492890472311C8E49251289248231140A05020140A04020140C4B29265C72AB7D",
            INIT_RAM_12 => X"AED56AB44A6556AB55AAD76CB65B2DB6DB6D6A37198C35DAED76BB5DACD66AB51A4CF46A",
            INIT_RAM_13 => X"AED569B45A251279349A4B2391475AC8F2793CA25129A5D3CE2996E7FDFFFFFFFF1B5D5D",
            INIT_RAM_14 => X"3CB0A396DC2E3B5DC7EBF3F6F9EC35FAFD6DB6DD6DB5DA6D32793CA2536BB65BF61B0D6D",
            INIT_RAM_15 => X"5DAED66AB499E8B2491C90472391C8E47239188E472391C8C45028100804028100C06041",
            INIT_RAM_16 => X"FFFDFFFCFD7536AB75AAD56AB4CAAD56AB55AED96CB65B2DB6DB6D6231186BB59ACD66BB",
            INIT_RAM_17 => X"A25129B5DC35FB0D96BAD569B45A24D269248E451C6AA409A4D27140A2554CA79E575DE7",
            INIT_RAM_18 => X"24944C271411C524DB9A5F70DAEE3F3F8FBED361AFD75B6DB6DB6DBADFB0D75BAD96893C",
            INIT_RAM_19 => X"6231176B359ACD66BB5DB0D66AB451C892391C8E472311C8C46231188C462391C9048241",
            INIT_RAM_1A => X"40A8964AABEEFBFFFFFFFBF4D8D9A4F29934A25369B55AAD76BB55AED76BB5DB2DB6DB75",
            INIT_RAM_1B => X"C365B3D9ED767AAB349E4F28955B6EFF4D86BF5769B3C9A4B2390471AA90271349A4E279",
            INIT_RAM_1C => X"2C9A4F4924D28954BA65B4DC6CB65BEE897DCB6FB9FC6D367B0D75BADD6EB6DBADF70D86",
            INIT_RAM_1D => X"AAD56CB65B2D96CB6D6631176BB59AED66BB6231186AB451A88231188C46231188C47241",
            INIT_RAM_1E => X"3C9A4D269349A4E271452A9E77DE7FFFFFFFDB6FA0724924D279349E5128944A25369B55",
            INIT_RAM_1F => X"BADF6FB7DBEDFB0D7DBEDFB0D96DB71F6D459A4B27945AEE5B9FDFDFE1A9B4596431B6AA",
            INIT_RAM_20 => X"188E48251309A504A25D34DD6FB824323924964B208FB9A5F73DC6E7EDB2D85BADD6DB6D",
            INIT_RAM_21 => X"9A4F28945A6D369B44AAD56AB5DAAD96DB6D6630D86C361AED86C36233176AB451648231",
            INIT_RAM_22 => X"F7F5E9B2C79AE9146934984D269349C5149240D332DDFFFFFFBFAE9640E17148E492492C",
            INIT_RAM_23 => X"C6DD6CB6DB6DB6EB6DB2D96BB65AAD1679349A4D28B55BEEDBBF759A4B2693CAAEBBDFEF",
            INIT_RAM_24 => X"6A33198AB491C8C2713D22944B261B6DE90C924D28B4DA6D36AB55AAC924965C76FB9FB6",
            INIT_RAM_25 => X"6DB6DD6F381C52392C964B259349E4F27934AAD16AB4DA6D56BB656633188C36631198CC",
            INIT_RAM_26 => X"9649239349E557EFD7F7F9EEADB491A4C26130984C2714526924B2B6F3FFFFFFBEDB6CC2",
            INIT_RAM_27 => X"8E4D2FBAEE3EFB1D75AED76CB75B6DB6BB55A6CD218E361A8924924D28964C371C125934",
            INIT_RAM_28 => X"6635198CC66351A8D46E371B8D365AED76CB71BCE0914924F69B5DB2D96DB6DB6D96CB4D",
            INIT_RAM_29 => X"F3FFFFFC6C6A4954B25D329B6E375BEE07148E4B24924924B2592C9E4F29B4DA2D36AB55",
            INIT_RAM_2A => X"349A4D2713CA2934B26134DC7038E4D36D96BB5FA686130984B2592C9C514A2512067996",
            INIT_RAM_2B => X"BB5FAED76BB5B6AB14A26377DCECF5F6CB5DAED76CB65AAD568B2C71AA8F269349A4D269",
            INIT_RAM_2C => X"8E4922924965129B556E371B8DC6A33198D4723F2291C8E472392C9ED36AB5DB2DD6ED76",
            INIT_RAM_2D => X"40A6944A240D576DE7FBF3F3D5540A49149A592C994C271BADF7038A45229148E4523914",
            INIT_RAM_2E => X"389A4C2592C964B2592C964B25930984C261309C4F2924D26944A2409A4C2592C964B261",
            INIT_RAM_2F => X"BADFB0D86C361B0D86BF5FAFD7EBF556394CCF73F8D96C2DB6CB65AED96DB5DA6CB1D6A2",
            INIT_RAM_30 => X"81BEDF6F371B8DA6DB65B2D84D36DBEE29346E371B8DC6E351A8D47A4769B5DAED76CB6D",
            INIT_RAM_31 => X"30964A25128944D28A512A934F3AAF5FFFF7E3594C2813CA0512894D28964C265B8DD6F3",
            INIT_RAM_32 => X"B6DF70D7D9230CF26130964B25128944A25128944A25128944925128944A25128964C261",
            INIT_RAM_33 => X"7E4D6CB86C761B1D8EC765B1D8EC761B0D7EC35FAFD76AECB2BBAEE7EFB1B7DBAD96CB6D",
            INIT_RAM_34 => X"4528944BA5936DB6EB6DB4D74AA55289449A4D269248940A2514B272371B8D46A351A8D4",
            INIT_RAM_35 => X"24924924924924A251289249249289A544A25122A699EF3FFF6D3C69A04F279409C50281",
            INIT_RAM_36 => X"DB636FB7DB6DB6EB7DC763ABB14551A4B25128944A249249248049249249249201248049",
            INIT_RAM_37 => X"6A33198D46633196CB7E516ED9ECF67B3D96CF65B2D8EBF5DAED76BF5FAFD55925B75DCF",
            INIT_RAM_38 => X"3C9E4E271389A4D2713CA0544B2592C996D3612A924813C9C4F279389E4F2793CA050289",
            INIT_RAM_39 => X"1C0E070381C0E080402010080401C100804920100804030A49349A555338DF7E7DF59481",
            INIT_RAM_3A => X"B75DAAB34AAEDB9FBECAE16FB75B6DD6FB96C7575E69234964A2512492480401C0E07038",
            INIT_RAM_3B => X"389C4F2793C9E4F2796E371B8D46A32D96CB7E4F6FD9ECF69B3D96CB63B1D86B7596BB65",
            INIT_RAM_3C => X"D377FFFB66DA0502793C9E4F271389A4D26938A05149A552C974C255228F261349A4E271",
            INIT_RAM_3D => X"2010080401C0E07038180C06030180C060301C0E08038180C070402010080493CB091513",
            INIT_RAM_3E => X"C763B0D76AED367B45AED366965D373F8DC6DB67B0B85BEE1B3D9EB2BCD14612C944A249",
            INIT_RAM_3F => X"449C4D261349A4C261349A4D269389E4E27976391C8DC6A32D86CB7E4F6FD9ED369B3D96"
        )
        port map (
            DO => promx9_inst_9_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => promx9_inst_9_AD_i
        );

    promx9_inst_10: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"2010080596122ADBC6FBFBE68813C9E4F2713C9C4E271349A4D261309C4D2794D2A954AA",
            INIT_RAM_01 => X"79A68D2592892492401C0E07038180C07030140C06028180C05028140C06030180E07038",
            INIT_RAM_02 => X"7E4F6FD9ED367B3D96C761AED65A2C72090482472ABA6EBF3B7DBEE36DB4DA6CF6BB5D65",
            INIT_RAM_03 => X"2C9C4E26938A25249A3C9A4B261309A4C26130984D269349A4D2717A3D1E8EC7237196C3",
            INIT_RAM_04 => X"140A06030140C06038201009261966BBCFFFDB3AD0279389C4D271389C4E279389E4D261",
            INIT_RAM_05 => X"DF71B8DAEDB6BAEB04511A4B2512490080401C0E07030180C06028140A05028140A04028",
            INIT_RAM_06 => X"823F1F8F476391A6C37E516FDA6D367B4D9EC75FACB458A3CDC6D37DD333DD7F3F3B8DBE",
            INIT_RAM_07 => X"389A4E269389A4E26930964C26130985027934984B2592C964C2592C964C26130964B261",
            INIT_RAM_08 => X"288E04020100804028140805028140C060381C1253585D77FFDF6549228F27130984D271",
            INIT_RAM_09 => X"9A5F77DDFEB6FB8DD6EB75B8DBEDB65A48B23C964A2512010070381C0E060302C9E4E269",
            INIT_RAM_0A => X"2C944B25128944A25182411F8FC7A391A8C3764F6ED96CF67B2D8EBF5967B0C75B8DA6E3",
            INIT_RAM_0B => X"409E4F269349A4E269309A4C261389A4D27138964C25928944D2592C944A25928984B259",
            INIT_RAM_0C => X"34BCE8955AED76AB54A24F248D23C9443020100A04020100806038203EF0BF7FFF39E681",
            INIT_RAM_0D => X"B6D1608DB69B4DA714BAE9BBFDEE371BADDEE771B9FE7CF4F5A692349449249201007038",
            INIT_RAM_0E => X"28944A2512C944A2592C944A25128144A2518AC3608FC7A391A6BB6DC92CB8ECB63B0D7E",
            INIT_RAM_0F => X"B2FBFEFF7CB2E8E271409C4C271349A4D269349A4B2592C9C4E27934944925128944A259",
            INIT_RAM_10 => X"2892480401C10185149E4D239148A472592C9647206FB85C0D7489288602018100A060D3",
            INIT_RAM_11 => X"65C52AB7EBB5B6BB4D9EC51B6D369B4DF755D375BBFCEE779FDFB6DB71B9FDFC73AD4471",
            INIT_RAM_12 => X"1C100904824924A25128944A24924924925128944A0482412090488AC5618FC7A37186AB",
            INIT_RAM_13 => X"61248C2401C2CB0BDFF7FFFFF143C964C269389C4C2592C964C261349A4704830964D269",
            INIT_RAM_14 => X"E7F5F9F968E2E9146124924804069C5259138A472593CA6532993479B092289449C554EB",
            INIT_RAM_15 => X"8AC762B047A34D66A259BF25B55AACF649248E49239148E452798EDF73B7DC6EB79F9DB6",
            INIT_RAM_16 => X"309A480591C184804020100804020120905124924A24824120924824164D2814C9C47038",
            INIT_RAM_17 => X"552A932994CA4502795542E595DCB65B8FE7FBEB9644024144B271389C4D2592C984C261",
            INIT_RAM_18 => X"DF69B4DAED765B9DD7EBF3F0D2465A48E25924901751C963CE1714964F2A954A2491E6BA",
            INIT_RAM_19 => X"54A8572D2652E572B18EC7629047630D569A5134E09359EC922924A2D56CB65AAD36DBAE",
            INIT_RAM_1A => X"30984C26128984C2592C984D2403096470381C0E070381C10090482410090513CA8542A9",
            INIT_RAM_1B => X"9A4F2490B79B0942AA50A6522994CA4512813896133138DD971B9EAE9E4704020144A261",
            INIT_RAM_1C => X"B6E3B1D8EBAD571DB6CF5D70B86B6E7BBFCFDB5B648E3551E4C2512CC7278F375BEE0714",
            INIT_RAM_1D => X"2012080894CAC542A954AA562B16D349C4DA8EC762B04722ED448A452A9D714964F28B55",
            INIT_RAM_1E => X"200C0603820120A2512C9A4C26128924C2512C984B240309A49030180C060381C1008040",
            INIT_RAM_1F => X"9E491D6F381C3216FB71B0974AA48A4532A148A2542A94CA04E27134980C0586540E890C",
            INIT_RAM_20 => X"452A9D724A6D76CB86CB67B2D8EB6D973D9EB6D970D75C371B8D9EA2C51F6CB4D1C4B2BA",
            INIT_RAM_21 => X"140C060381C0E07038200E142B95CAA572CA60B0592C1793A9D4FA96C963B0C762ED3482",
            INIT_RAM_22 => X"40960B050202E9A430100A060281C12090482C984C25924924A2612C964D2914CA651279",
            INIT_RAM_23 => X"8E411C6B2491A6174475B8DD6FB81B8D649144A25128944A2512DAAA6570B5C9DC6DD4A9",
            INIT_RAM_24 => X"9ACB64B0C7630D24A265BEE4945AEDB6FD8ECB65B3D75AADB71D86AAD36BB86DB69AFB3C",
            INIT_RAM_25 => X"2C1C152A950AA93281388805030180C07038142A532B960AE582DA71369A4F281429F513",
            INIT_RAM_26 => X"DF6FB5B8DB650E570264AA4E040200E112200C06040281C120904024184C24928944A251",
            INIT_RAM_27 => X"A6D36DBBECB5767914863EDA6A240C9288D379BEDF6E355204F279389C4F28140A86DBBE",
            INIT_RAM_28 => X"813EA15028544A57239ECF66B257E34D76DB824B2AB65BADB6DB75C767B3D65AADF70D6D",
            INIT_RAM_29 => X"24164B26130944A0483024564BA592C95299489E44028180A070794CA6572C164B29D4FA",
            INIT_RAM_2A => X"389C4D271595D76DA5DB6770B75A650E571B793C95270201208030080603020201208040",
            INIT_RAM_2B => X"C765B2D75AADF6FB5DA2D973D85AACD2290C823AD96A29A4F1B6F379BCD9491389C4E271",
            INIT_RAM_2C => X"60B0592E26D38A15028DCAE67338D48E673BA2D167B2D8A3D1D90496556DB75BADB6ED86",
            INIT_RAM_2D => X"0C060202018100804020144B25128940708950AA974BA612C964AA4CA44F228140A102A9",
            INIT_RAM_2E => X"6DAC8F271349A4D26930984B0DAB66572B85BE616E96CAA50E57238540962883C1207050",
            INIT_RAM_2F => X"9A556CB7DC361B0D8ECB69B2D6DAADB6CB45AADD6CB3C96472290C7DBAD973C9A38DD6FB",
            INIT_RAM_30 => X"50A651271102C5B4C15CAA5C5028146E573395CCE6733AA532B954A2D369B3D96C72391C",
            INIT_RAM_31 => X"793E9C491489A07038100402018140E0804020100804828921029954B0994CA6130974BA",
            INIT_RAM_32 => X"7DB6E893C71BCDE6E3551C4D27134984C2582C141855CB25D2D97CBE5B2B95CAA50E6723",
            INIT_RAM_33 => X"AAD56AB459ECD66B45A6D76EB8ECF67B3D9ECF6BB2D65AAD56BB4DAAD36592C924521904",
            INIT_RAM_34 => X"61329A4D2692E984B254A65127165369C4D168BEA472B95D2E7733AA50EA954AE572C95C",
            INIT_RAM_35 => X"B254EA75CAA55267438D429D4A950A00C0301C0402018100E070401C1008048201E542BA",
            INIT_RAM_36 => X"AACB2492C8E452290C79D1288EB79C0DD6B2409C4D26130984B0582C166675C81CEEB97C",
            INIT_RAM_37 => X"A6552D975BA5D6D96CAAD569B45A6D56BB65B6DD71D96CF67B3D9ECF69B2D5DAAD36BB6D",
            INIT_RAM_38 => X"180E070583C2A584CA69349C4D26934994C259284E1028DC09C4F291C4A253391D52E944",
            INIT_RAM_39 => X"28246A96C79C0E876CA9D72E985C6E16C94395C4E66B95CA250248180402018100A06038",
            INIT_RAM_3A => X"D369B0D5DA6D36AB4DA2492491C8E45218FB9E531C6FB81BED8491389A4D2592C160B050",
            INIT_RAM_3B => X"8948DF51B99D0E796CAA572DB7DBEE56EB85AACF6693DA6DB6FD86C761B1D96CB65B3D9E",
            INIT_RAM_3C => X"1C0202018100A060381C100A0894CAC584C269349B4DA6D34994C259266051399C6E472B",
            INIT_RAM_3D => X"349A4C2582C140A05024246676481BCE275CB2572C96CBA5B2C9649DC4E04E25CAA51281",
            INIT_RAM_3E => X"CB63B1D8EC765B3D9ED367AFB55A6CF269248E472391C8E452192CA240DF70B81BAD7481",
            INIT_RAM_3F => X"594AE8764A64AE671B95C2A151B9DCEE8954AA6172B95CADF6DB75AACB22924A2DD71D96"
        )
        port map (
            DO => promx9_inst_10_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_5,
            RESET => reset,
            AD => promx9_inst_10_AD_i
        );

    promx9_inst_11: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"A5CAE14EA6D30542912C0202018100A060382024522A950B09A4C265349B4DA6D36994C2",
            INIT_RAM_01 => X"9A40E27137DB8D5471349A4C2602C160A0502424637236D329C53BA1D2F1995A5CCEA95C",
            INIT_RAM_02 => X"AAC9209149AD96FD8EC761B0D8EC767B3DA6CF67AEB55A247229148A472391C8A432193C",
            INIT_RAM_03 => X"69349B4E2713ADA4BA4CCAE8944A6552872B91C6E472395CF2794C924D29985BAE574D8D",
            INIT_RAM_04 => X"754AEA74BA9D0E875CA1CCE46FA713495291340402018140C060504CAC5A4BA5D28964CA",
            INIT_RAM_05 => X"8A452391C8E432793C85C6E491B85BAD4479389A4C0582C180B048281E5D51B68AA58302",
            INIT_RAM_06 => X"8A34EFB6DAA5F72B85AECD609048A516DB86C35FAFD86C765B3D96CB63AEB4C9A4721914",
            INIT_RAM_07 => X"50AE574B25D26584CA69329C4E275B8994BA48C8E89548DD52893C99C0A1723A6531D575",
            INIT_RAM_08 => X"3012112D26120562F27D3EA4543AE592A95CB24AE470A7936962993C8202018140A06078",
            INIT_RAM_09 => X"BF5DAAB449A432070C8A45229148A4D2991B8DC92592489BAD54914CA85329950AA55291",
            INIT_RAM_0A => X"9DCAE573CB2552073C7A2AAED1BB6552DB75AED1618F3824D2CB76C35FAFD86C765B1D86",
            INIT_RAM_0B => X"380202018100C1227058AC564BA6130984CA65349B4E26930984B250CD2893C9E512673C",
            INIT_RAM_0C => X"793A9C4DA6934984B24C9A090A9652CD72C968B8A2564B6592C964AA4EE571B7D3497299",
            INIT_RAM_0D => X"BF5B6CB6DBB61B0D7EBF5968B3C923EDF70C86452190C865328913924B2592C8DC4DF4FA",
            INIT_RAM_0E => X"4CA05F7349E4B2572399C6E672B9E4ADA449619652564B25B6A95CAED1628F37E4B2AB76",
            INIT_RAM_0F => X"9DD0E872385B897299340402018101A122A150AC984BA5D2E984C26932994CA653095299",
            INIT_RAM_10 => X"9A4F2893C99C8E2703813C9E4E26D36994B9549C46089552A952C954AE61533BE5D2775C",
            INIT_RAM_11 => X"AACF618EB79C528B55B2D76AB65B6DFB0D7EBF5768B3C9240DF7038643207039E5323724",
            INIT_RAM_12 => X"6132994BA5D2A53299409E4810391C4E472B91CCE37236D46E672B5D228B313AE4B2794C",
            INIT_RAM_13 => X"5938E5754A1E371B7DA1D0E671B81B6952892004040202422542A154AC984BA6130984C2",
            INIT_RAM_14 => X"8A40E06FBA2512272CAA596DB4C99C8E371385BE9E4F275369A4BA58A44806054AA5B4F2",
            INIT_RAM_15 => X"5D104D313AA53279239EC91E6D36DC126B5DB2D76BB65BAE1B1D8EBB4F259449A4522914",
            INIT_RAM_16 => X"612C964BA612E984B26132974B254A647028349A010007DB8A471B85C4E271391C6E2713",
            INIT_RAM_17 => X"5CAA4D25040AA5B4FA613ADB71B81B8A4733A1C8E46EA652C512600C06030282C26542A1",
            INIT_RAM_18 => X"9A452593C96492592C92472192CA242E373CAA5B6DB4C9DC8E471389C2E06FA793A9B4CA",
            INIT_RAM_19 => X"7D42E070B81C2E27138D926070375C2E27039EC91D6CB6DBF27B5DB6DB6CB76C363B0D6D",
            INIT_RAM_1A => X"0806050281828564A94CAA552A95D2E974B2612A552A94CA2450381004030180038A16F2",
            INIT_RAM_1B => X"8DC6E271381BE9D4DA60A84D2603424552B960BCDA4EA9E552992B8138972B14CA24C020",
            INIT_RAM_1C => X"C361AED76BF5B68B0C81C9259148A472592C9A4B2394CA242E4944AE5B6C94CA1CEE6723",
            INIT_RAM_1D => X"180600000000E1B4F2713E9D5037D3E9F50381A85F7037DB89D4D29ECB1F8DB6DC128B6D",
            INIT_RAM_1E => X"5CA853291409402010100A060381828552B254AA552A954AA562A954AA5329944A044030",
            INIT_RAM_1F => X"AE596B954AA50E893B95CAE471B85BC9D4DA652C532802C140C08144A6562B160B29B4C1",
            INIT_RAM_20 => X"A6D1638FC79C528B75BF61AEB6DAEC91F70B8A43206FB81C52392C964B259559A44E594C",
            INIT_RAM_21 => X"50A65228940960A06030225129144A04F2B269369A4DA6D389C4EA71369C4E2713697280",
            INIT_RAM_22 => X"2C180D07044A65229148A2502681C02010180C0E142994CA0542A950A8542A954AA552A9",
            INIT_RAM_23 => X"92492795585C6E6954B6DB6C96CAE552A94C9DCCE572389BE9D4DA652C54289300E07048",
            INIT_RAM_24 => X"6D369B4CA6126552B1A6D3658FC7DC52796DC361ADB458A3CE170B7DBEDF6FB864523924",
            INIT_RAM_25 => X"7538972A150A65329148A4512792C1E4F2894CAA5528148A85429944AC562B96930994D2",
            INIT_RAM_26 => X"64AC54289340E0603020140B068381E0F07038180A0380800010B17146C710391C4DE4FA",
            INIT_RAM_27 => X"7DBEE070C86432291C8E4728B4C7DC6E7954B2D72B96CB2552A94C9DCAE471B85BC9D4D2",
            INIT_RAM_28 => X"50A8522A154B48E0CA6534974304CA6542B1AAD3648FC79C327B65BF5DA7AFB79C0E06FB",
            INIT_RAM_29 => X"85080D27195C6E2702813A9D4C954A452289449E4E25038A25329954A8562A94CA8552A1",
            INIT_RAM_2A => X"91C8E2713813C9B4D260AC53281301006030180C070402814090401C0A0601800226350A",
            INIT_RAM_2B => X"B6D5606F381BEDE6FB81C0E170B81C32190C8A432793C75C4E5954B2D72B974B2572A943",
            INIT_RAM_2C => X"54A8542A950A6552A94CA65329150A2512702816070A154AA52291AAD3648FB79C326965",
            INIT_RAM_2D => X"2010030A995C8E4681511A6571B91CAE271B81429E4E264A25027930180A0793CA253299",
            INIT_RAM_2E => X"B6DB6D96CAE52EA7338DC6E2713813C9C4CA60AC532782C0C05028140C06030140C07038",
            INIT_RAM_2F => X"B2D5659047E4125945A6C51E6FB79BCDE70385C2E170381C0E070C8640E692C75C2E6954",
            INIT_RAM_30 => X"18140D0793C205229950A6532A14CA8562A150A8532A150A451289381E542A93C9E562D1",
            INIT_RAM_31 => X"140C0B0713CA050281382A6570A91CEE56DB34A2A573395CCE471B85C49E4E26D3049048",
            INIT_RAM_32 => X"81BEE69246D40E493CA2532B96CAA4EE973B91C4A04FA793C9C4D260AC51268300E05028",
            INIT_RAM_33 => X"3C20562B160AE5B4E2BF5967B14824323924863EE06F37DBEE070B85C0DF70381C0E0703",
            INIT_RAM_34 => X"89C4E04F26D349822814160C070341E0E0893C245229148A8522A94CA45329150A653299",
            INIT_RAM_35 => X"50AA51280300E040201C164D2914CA4522DA794EEE95CA5D2E774B95D4E873B9DD0E7733",
            INIT_RAM_36 => X"81C0DF6FB7DBEDF6FB7DBCE7924653CE172492492896CA5C6A67338DBE9F4EA71389B4A9",
            INIT_RAM_37 => X"4CAC5729144A45128954AE5A47058B25D4F2C35B68B248243219047DC31F6F37DC0E0703",
            INIT_RAM_38 => X"AE572A94CA5D0E874395C2E370A7534982890C140B068301E0E0894022500684CA452289",
            INIT_RAM_39 => X"853C9D4EA6D349A4B154AA522803412040383C9E5026954AA614C995D2E9733ADD52C954",
            INIT_RAM_3A => X"8E42DF6FB81C0E07037DBEDF6FB7DBEDE6FB7DBEE592465369D70381C0E5764AA4AE6723",
            INIT_RAM_3B => X"40A2100783426562C15CB25A4E254A2512895CB4972DA713C8D312C35B68B2C82411F904",
            INIT_RAM_3C => X"79572C974B65F2D95CB65B2D964AE572994BA1CCE3723853C9A4B9101607050301E0F078",
            INIT_RAM_3D => X"79BCE275CA650E8723853E9D4DA6D34994C158AA5327830120B0814CA8542B2653EA673B",
            INIT_RAM_3E => X"BF5969B2C863EDF9148E40DF6FB81C0E06FB7DBEDF6F37DBCDE6FB7DBEE493C69309A4E3",
            INIT_RAM_3F => X"20120B0402C1A0C060381C0F0A15CB4992C160AE5A4EA7130532A964B69E4D17D42A1522"
        )
        port map (
            DO => promx9_inst_11_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_7,
            RESET => reset,
            AD => promx9_inst_11_AD_i
        );

    promx9_inst_12: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"48AA9A4D2654CEA76CB65B2E964C66132B5450DD2D974B6592C95CAA50E672B89BE9C4B1",
            INIT_RAM_01 => X"79BCE074C922E984D271BADE744A5CAE57127D3A9A4C964B2594C158A852280301C152B2",
            INIT_RAM_02 => X"60C29B4B96D4AE574BBF5B6AB348A3CE19248A3EDD6F381C0DF6FB79BCDE6F379BCDE6F3",
            INIT_RAM_03 => X"B654E873B91C09C4C920120B03828180D068342A542B9509C5A4D1793A9C4EA75389B4B1",
            INIT_RAM_04 => X"58A652280342C594D2712C9A4F2A5D93097CA66B71B84CEDF34B5CCEE12F96CB65D2E974",
            INIT_RAM_05 => X"79BCDE6EB79BCDD6EB75B8DC7349A30974C2653099523A1C8E47127D38992B958AC562B9",
            INIT_RAM_06 => X"7940A272B813C9C4A928964F28A8554ED974BB5B6BB3D8E3CE392485BADC6F381C0E06F3",
            INIT_RAM_07 => X"BE6775B95BE612F97CB6592B94399C29F4DA28120A03820160D0A94CAA5C4B94CBA8E271",
            INIT_RAM_08 => X"7936582B14CA6552A954A6522804CB09B4EA793EE074C8DE572B6D65E573B9DDAE972BB5",
            INIT_RAM_09 => X"7DB8DC6F381C0DF6F379BCDD6EB75BADC6E36DB8DC6FB9E49164B2592A964EB99C6E570A",
            INIT_RAM_0A => X"4CB0562A97946C92B260CAE671389C4CB0E22C944F33BA1DD3399CB7596BB3C8E3CE3924",
            INIT_RAM_0B => X"A2D135BADD6EDB5B34926775BA5CEE130984BA5D2D94B99C6E04EA28140A0582026510A9",
            INIT_RAM_0C => X"5D2E944BA89C4E24EA7534972B954A6552A150A45008954B09B4F37DC4E4754BEDF74BA5",
            INIT_RAM_0D => X"B6D96BB3D8A3EE492C7DBADC6F37DBEDE6F375BADD6EB75B8DB6DB71B8DC6DB8E51268BA",
            INIT_RAM_0E => X"24120904054A4162B158B05D4E2854ADC53B95CCE774399CEE572B713896343B65F319A5",
            INIT_RAM_0F => X"81C2E897DCEDD73BADE777B6DC6DB6B77DEF766977B859DE773B95C2DF2E964A5CCE0448",
            INIT_RAM_10 => X"71B8DB6DB65C72792C89B494491613EA04EA6D34992B958A8552A14CA00F09150AE9C4F2",
            INIT_RAM_11 => X"A1C6A6753856377BA5B6D76BB3D8A3EE49247DB8DC6F37DBEDE6F375BADD6EB71B4DB6DB",
            INIT_RAM_12 => X"CEE371B74B24ADD4382814090A154AA552F264C09C523794AE6753A1D0E8754AA52E7743",
            INIT_RAM_13 => X"44200F091592C9B4EA85C0E794CC6E772BB6DF6DB6DBED2FDF6C50C26D77BADE36973B9D",
            INIT_RAM_14 => X"75BADD6E371B6DB6DB6DB6DB6D365B2DC70B81C2DB6994CB29E4E26D349A4C158AA54299",
            INIT_RAM_15 => X"65572C95CAA5929754AE52E977CCAE776BDEB2D76AB3C8E3CE492C7DB6DB6EB79BCDD6EB",
            INIT_RAM_16 => X"E36FB4B9DDAEB75BADDAE974B8CC644962482812182B154AA5C4898D48E471B99D327651",
            INIT_RAM_17 => X"6D34982B958AA5429148A00D08958B09B4FA85C6E572BBA675E57DD2E775DBEDB6B77D3B",
            INIT_RAM_18 => X"7DB6DA6E375BCDD6EB71BADC6E371B6DA6DB6DB6DB6D365B0D74AA5538D94A144A65B4E2",
            INIT_RAM_19 => X"454CD0261A1D2E976CA2164418CBA592E96CB65929784CEED7ADB5B2D56AB34923EE492C",
            INIT_RAM_1A => X"BAE579DCEDF71B6DC6E777EB9F7DB6776DB6D6E773B9D8534480482428582D14C3AA76AA",
            INIT_RAM_1B => X"492C9A4C248A4572D26D32572B154A85228940980908954AA584DA81C2E174495D51F77D",
            INIT_RAM_1C => X"AED56AB3D923EE292C81B6D96DB75BADC6DB71B6DB6DB69B4DA6D369B4DA6CB6130964A2",
            INIT_RAM_1D => X"1C30614F26CBEA349279D72991BAE5B2976CB2676E984C6DF2D964BA5B2977CD2ED77BB5",
            INIT_RAM_1E => X"79C2E472385C6ED923CAE975B9DDF6DB3BE7E3656E9BEE76375B85DAEFB2B12509409048",
            INIT_RAM_1F => X"65B2D96C25D2C9549A55389F6EA6934984C164B0562A950A65228138180B07954AA552DA",
            INIT_RAM_20 => X"B6592B743BE6F76BC6B2D76BB4D963F2072C8636D84C26DB8DB6D369B4D96C26130994CB",
            INIT_RAM_21 => X"D6E51D46034120A050693EA24FA954ED755B6D5B2A964B2572977CBA5F34B7CBE6971B84",
            INIT_RAM_22 => X"3C9A0C07050A6532A1653AA274C8DC4E376C95DF6FBA6C2F1B9DEFFFF9F4B9DDB75B9DA5",
            INIT_RAM_23 => X"6130984C25D2E984C26530984BA592A9449A6D44E26FA75389A4C15CAC552A948A451281",
            INIT_RAM_24 => X"CAE371B9DC2DD6D954BE6132860AE4AF6B9DB3596CB4D9E411F7248E38D74B26134D96C2",
            INIT_RAM_25 => X"BEEFB6B8DCAEB6E9849D9E142B960AC54258894AA253B91BCF5B64C65B2D96CC20E32B43",
            INIT_RAM_26 => X"652E572A950A652289409C4D07048A65228148AE9B4FB75A8912DAAE512A95CB65733B95",
            INIT_RAM_27 => X"923ED74AA5930974B2592C974BA5D2C974B25D2C964AA5528924BA89CCE571B813C9C4D2",
            INIT_RAM_28 => X"BE552376C9DDB38D95D2E773B8DCAE76E93CC2592F838404AF5BBEAED76CB559EC51F71C",
            INIT_RAM_29 => X"38BAAA943A24EE995CBE5B2B94B9DC69D4B15CB25A4EA6D32582B1894CE773BA5BAE377C",
            INIT_RAM_2A => X"A2512772B8DC09D4E26932972B150A853289409E4E0683CA4512703CA2532A9549C4E268",
            INIT_RAM_2B => X"AED76BB55A2C71E7048E42D96AA552C954AA552A954AA552A954AA592C954A24D24924EB",
            INIT_RAM_2C => X"A1D2EC753915B289ADCAB8E48B3AE6966995DAE97AD9DCEE1309BDBE5B1C499549C121AD",
            INIT_RAM_2D => X"382451289449C0E0601C120A0388146E24FA853C9E4EA58A85B4EA64BEA0502813A9B4C9",
            INIT_RAM_2E => X"51289349A492292513AA532873391C29E4E26932982B154A85329144A04E068341E10080",
            INIT_RAM_2F => X"BE52D20A958AE592D1B2D76AB4D9EC71E6F386451C6B2512A954A25128944A25128944A2",
            INIT_RAM_30 => X"8DC8E271295C29B4D1CE52EC75BC25F31B54DEC91C6FCD6E7607C6DEEB74B8DD2E56A995",
            INIT_RAM_31 => X"44A04E06830180E07838180E0702C140803024140F2793CA04F2683414070A160BC9E512",
            INIT_RAM_32 => X"5128944A24D269349A4D269349145205132BB6572A94395C4A04EA6D32982B154A854291",
            INIT_RAM_33 => X"DF6B73B85C25B2E99DBA54D42B960B69D4E2B7596AB4D9E491E6EB86451F6C25126944A2",
            INIT_RAM_34 => X"389C142C16D42A272395C8E36E291C09F4EABA4EE673BB644B4BBDDB3F2BBDEC6F5B6B2B",
            INIT_RAM_35 => X"6932562B154A853289409C0E0602C120A0683C1E0D060240C0504034A2522894CA04C081",
            INIT_RAM_36 => X"7DC5228E35528934A2512A944A25126944A251269348A45205153CC2DB2B95391C29E4E2",
            INIT_RAM_37 => X"CEE377D95D6F3B6DADD6ED71BBDDB6976B6C6CD4D72C168B25E502BB5BAAB4D9EC91F8EB",
            INIT_RAM_38 => X"50961029150A65229144A0552D27946E670B95C8E472391C6E04FAB1DD35BA5ADEB79DBE",
            INIT_RAM_39 => X"C2D3132D2713A9F4EA75389B4D164AE542994496090502C0C03050341A0D0581C0E0C089",
            INIT_RAM_3A => X"BF5DACB4D9E471F6EB7DC5238FB612A944AA552A954AA552A954AA552A94492492051334",
            INIT_RAM_3B => X"CE6135BADDF7177DB5CEE776DC6CAD534BD6D6F7AF9B5DF6772B7CBA52C80C96CBC9F502",
            INIT_RAM_3C => X"28180C0602C16152A950AA552A954A85329148A2562C97D46E67339DCAE572391C8E14E2",
            INIT_RAM_3D => X"592A944A24922522F385284A261613EA05027D389C4D968AE502914CA44F05828120A050",
            INIT_RAM_3E => X"B638992DA7540A151ABF5FACB559EC71E6E379C0E16F3652A954B2592E964BA5D2E974B2",
            INIT_RAM_3F => X"9DCAE573391CAE36DADEE974B84DAE976D54EF73AB985C6F7B6BADE36FB4BB5DAE571AFB"
        )
        port map (
            DO => promx9_inst_12_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_9,
            RESET => reset,
            AD => promx9_inst_12_AD_i
        );

    promx9_inst_13: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"48A855299449A0B0602C140A0502420542A950AC974B158AC5029944A6582DA8548E874C",
            INIT_RAM_01 => X"5D2E974BA592C964B2552A9449A453CD426930AC974386D44E05127D3A9F4F260B49B4CA",
            INIT_RAM_02 => X"DF71B6B8D6534F2B54AA2A5C4C9853CA251ABF61ADB559EC71E6E36DB6DB6D35D2A964B2",
            INIT_RAM_03 => X"4CAC5A4FA85C8E774C9DCCF6B4395CAE46FADEEB79DADE771B5B3CE37FF1BDEBEE579D95",
            INIT_RAM_04 => X"89365B4EA89409F4EA7136992B950A44E06030160B050302A552B1612E564B158AA552A1",
            INIT_RAM_05 => X"5D30984BA552A954B2592C964AA552A944A2512692492A1CEDA4BA95CCE572348C2D7512",
            INIT_RAM_06 => X"E36DB5B95EFEBBADAEDB6B75BDEBEE56F974A1B25E4FA8940A24EABF5FADD55A6CB1F6D3",
            INIT_RAM_07 => X"753C9425848AE552994CAE5A2F289CCE894CA6532A943A24AE47028DEB7FFDEDF6B71BE7",
            INIT_RAM_08 => X"9DCEE873B9DB8A573B95CEE673395C8E370A7D3C9C4D25CA85226838180C05844A855313",
            INIT_RAM_09 => X"BF5FADB559EC91E6BA592C974AA552A954AA5528944A251269349A49249134CB25728743",
            INIT_RAM_0A => X"30E574DBEE3617DFE7F7DB3BDD6D76976DCED2E973BBED2E76D94C7532563028944A571B",
            INIT_RAM_0B => X"38180C06850B4A36FA5D46E471B79305629850AC5B4EA91D729985B65B1454CA23CE1679",
            INIT_RAM_0C => X"49205E78CBE592A94BAE552A91B79D2E974BA1D0E8743A1CEE67238D409E4E260AC53280",
            INIT_RAM_0D => X"6D3A9F502754AE9723BF5FADD55A2C91C6AA552A954AA552A944A251269349A492692492",
            INIT_RAM_0E => X"B2591556C4D590927930E573B9DD779F3DCEE36FBEFCEE75D3ADB5E76572B85B6592A902",
            INIT_RAM_0F => X"8DC4A04F26D2E55289381C0C07854BCA171B8DC8E271B81C09A2B14CA85B4EA8DD0EA984",
            INIT_RAM_10 => X"492492492492291489409E74B95CEDB2B96CB65B28882A6592C953AE5715553A5D2E772B",
            INIT_RAM_11 => X"DAE173B5CC2D3276B969265E51399C2A5754BB5FAEB559EC71A69A5128944AA55289349A",
            INIT_RAM_12 => X"5CAC592E285CCF0B8DBEE99B74CB22249281140232BAEDF6DB9DBEDB6576DCEE36DB4BC6",
            INIT_RAM_13 => X"B24CE575BA9D0E772299C8E25026D3256289341C0E0818DCAD65238DC6E271B89C4E04E2",
            INIT_RAM_14 => X"4D26944AA51269249249229148940A0502793C9C74BAD89B4AA974BE5B1A492BA5D2F964",
            INIT_RAM_15 => X"C6EDAD985D2DD2E954B65F74B549DD0D92B96D20615239DD32672BB75DAED65A2C1154A2",
            INIT_RAM_16 => X"95C8E271391C6E3702792E582E285C8E99AEBAF5ACB6C593F1E8F4CB1E99585DB6BBBF9D",
            INIT_RAM_17 => X"6DAA8C2E3C6E32A984C25D2C964B1D4E773B9DCAE14F26CB056281381E0F3029DA88C313",
            INIT_RAM_18 => X"B75DAED75A2B4D349A4D289449A4D249148940A0502813C9E4F279349C6DBAD75A69D6BA",
            INIT_RAM_19 => X"8643144EBBEE379DBEB2572B93BA644E7744A1DF1F53B919A102A158BAA052B91CAE068A",
            INIT_RAM_1A => X"3C1E1F4E29DCCE773B99CAE57238DC8E3713813A972B138C8E79AEB2E16C91349572B923",
            INIT_RAM_1B => X"389A585ADA636DC8C3BEE77DFADD2E973B95CA612F96BB1D6EA74399C8A04EA713255278",
            INIT_RAM_1C => X"60B69B4F2AE4ED0386B2DBAED6D962A934924D269349A4922902813C9E4F2793C9C4E271",
            INIT_RAM_1D => X"D769B093485CEE77037D24524B2085929964A5D0E674391CECB12389C4D532B441A0C0A9",
            INIT_RAM_1E => X"A1CA9E4E268AE542784048D24CA99CEE89339DC6E572395CAE57238DC6DE4692CAC9F523",
            INIT_RAM_1F => X"3C9E4F271389A4E269349A513C6D6C522965D6F3B8DB5CEEB75B9DCEE331973ADD2A9753",
            INIT_RAM_20 => X"85C2D4268301A0C09958A8594EA8DBAA298EB2DBAED5D7DA492492492693492452050281",
            INIT_RAM_21 => X"95CAC90DA249E5C754CAF5ED97CB263637655D1E544791C161232B95CCE472391B6A571B",
            INIT_RAM_22 => X"DEF5B3984B1DAEC763A1C6A04E264AE520914032944EA95B8E573B99CCE673B99CEE7733",
            INIT_RAM_23 => X"49249248940A04F2793C9E4E271389C4D26934984C303DF71B8DBEE371B7DC6E76D78DA5",
            INIT_RAM_24 => X"301C172FA793C9E4B12C180E07038180C0704CAC572BA48B6A072CB75BADD4565A691492",
            INIT_RAM_25 => X"99CCE874BA1D528743A1CEE56EA48901E77DAAFFFBD3BA246D549A3CB09429948980C058",
            INIT_RAM_26 => X"DF77B9DEFE373B5BD6DEED74B9CC25CEA7539D449F4E168AC522914440DC70A99B49E523",
            INIT_RAM_27 => X"B75DADB2C552691492492491281409E4F2793C9E4E271349A4C26130964A29AE771BCDD6",
            INIT_RAM_28 => X"4CAC53291341A0D06834160D0602C1E0D068381C0E0783C200D068509A152B9652696503",
            INIT_RAM_29 => X"48AC5D72A79184E261A5CCD055CAA552B95CAE552973B8140A474CEFD55F72B719C59489",
            INIT_RAM_2A => X"30964A289D6F5B6DC6EB79BBDE7E76D75BBDD6E974984C258EA74B95409E4D964AA54291",
            INIT_RAM_2B => X"4CAC532B1651A512B2BB5DACB145124902894522912813C9E4F271389C4E26934984C261",
            INIT_RAM_2C => X"965F8C259209A4F2B958AA542782C38A15138944A05027D284E060381C0D070449E0D068",
            INIT_RAM_2D => X"8D409D4D964AC572B158AC6AB43390A0824138946F95CBA44EC974B6572E850203461764",
            INIT_RAM_2E => X"389C4D26934984C2592C964A279A273B8DDEF7F9BADE7F7F5B7BDED26330973B9D6EC73B",
            INIT_RAM_2F => X"6D220E07840A04E0803824522A958B2994CABF5FACB0451224F28140A0502793C9E4F271",
            INIT_RAM_30 => X"BE5F2E95CA1B8890D29E34E4AE365A04E0703820101137D2A5E50248C49F4FA7D3C9D4D2",
            INIT_RAM_31 => X"D6E733963B5DAEA73A95429F4E168B2592B95CA8696995DB2CA2926DB8E277CB24EEE974",
            INIT_RAM_32 => X"3C9E502793C9E4E271389A4D26130984C2592C944A2695D6778DE7EFFBB4BD6E37178DAD",
            INIT_RAM_33 => X"38AA5E4FA5CBC9D4F2793A992703C2251270301E112A154AE562E2C361ACB0451204F279",
            INIT_RAM_34 => X"7DD931B74CAE572B8DB66571B74AE4ACA078401E0C0783C1C10060402A5D4C144389A29A",
            INIT_RAM_35 => X"D6FDFDDE7EF75BADC5D6E92F77BB9E32774399C49C2D95CB0582C15CB2AA70AA122A18D2",
            INIT_RAM_36 => X"C763ADD0451224F2793C9C4E2793C9E4E271389A4D26130984B25928944925048B8AC9D6",
            INIT_RAM_37 => X"5CC4D72D968B89A2D96D345C4C960BC9F4FA7D389B4D244A251289401E0E0814CAA4E0B1",
            INIT_RAM_38 => X"64AC6B752994B08164CAE574B7CDAE9616CB69EB73B8DB646880803C20100803C1C0F080",
            INIT_RAM_39 => X"28924904038AE5D544EB79FEFC6F371BBDCEDEE72E76BB5D6EC753852A582B954AC5B2C9",
            INIT_RAM_3A => X"40A04F060401E132A1C361AED14512490281409E4E271389C4D269349A4D26130964B259",
            INIT_RAM_3B => X"402011080442211060893CA04C168B89C4F275389A2D16D3A9F4F27D3E9C4C96D2452260",
            INIT_RAM_3C => X"60B4592B154B05A2C964B257352C1D8EA994CEED75BDEAA696FBA5D6DF32BA5BA4AC8078",
            INIT_RAM_3D => X"34984C2612C964A25124920804028225A50295E77BDCEEB6FB7BC6E2E531974BA5AED91A",
            INIT_RAM_3E => X"793E9E4E271245129148A6500783C1C10088C363AED2C55228F2793C9E4E271389C4D269",
            INIT_RAM_3F => X"D6ED76B8DAE50C907840200F08044A21114B893A9E4C97538992EA75345A2D1713C9C4FA"
        )
        port map (
            DO => promx9_inst_13_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_11,
            RESET => reset,
            AD => promx9_inst_13_AD_i
        );

    promx9_inst_14: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"D6E12E9638DD92351A8534592C15CB25A2C964B25518CC654B39BDE2EF79DEEE3697CFAD",
            INIT_RAM_01 => X"389C4F269349A4D26930984B2592894492492412090482416132D27D369659DE371B6BDE",
            INIT_RAM_02 => X"70B6562C97D3A9E4F2793E9F4FA6D1C5429148A45128848AA562C1BF61AED4561248E269",
            INIT_RAM_03 => X"DF6B7BDCEF36F76B6DC35131B84B22C430703C224F088381C1113B7D2E5B2EA753A5C4E2",
            INIT_RAM_04 => X"6938984DA7548F0B8DCEE12B74BA1C6A872B8D385B2D164B0582E170B85734AC5EB38BA4",
            INIT_RAM_05 => X"BB5FAFD5D71A68E261349A4E26930984C26130984B2592C940A26144A2522994CA4532B1",
            INIT_RAM_06 => X"68BA604D98114080A96CB2552B164BC9F4E17540A1502813A8709948A0132A95CAE5C4EA",
            INIT_RAM_07 => X"74B05733AB5E339DC5D2F5B7DC6EF71BBFBEE375B4B84958C05068381E0F078401E2F933",
            INIT_RAM_08 => X"6130994CA6530584D275409A4DA813C9D4FA7D3E9E4D95CD7297438D3A5E4D970BA5B2C9",
            INIT_RAM_09 => X"3C2A5A2C160BC942D2BB5FB0D6D92268F269349A4D26130964C26130964B25930A0532B9",
            INIT_RAM_0A => X"44200E07840202F90A64C2A55126D264A28158B0562C15CAC5A2D98142A150A85368A089",
            INIT_RAM_0B => X"91409C2E96CBC9F4FA74B8582F1C5E0F199CDAF7B4BB5DF73BBDB5EF6FB3B5C7D389A268",
            INIT_RAM_0C => X"2C964B28154B29A4DA6D389B4DA6D369B4DA7544A34E28946A35127D3C9D4E16CDB28743",
            INIT_RAM_0D => X"7D3EA151A8D3E8E2705CB45C2B934984B2A1B75BB0D7EAAAE9026930984C2612C964C261",
            INIT_RAM_0E => X"E36B72B12893C9D4E26D30582A94898297028140A552A7D3C5350B34B05207868BA9C2FA",
            INIT_RAM_0F => X"81409A2E28DDB2972B913E9C3028D386150A74BEA050A855CF27A4E2F9BFFC6D76FB8DB6",
            INIT_RAM_10 => X"2C984C25930984C2593096532CA753C9E4FA7D3E9E4F271389E4F28546E47138DC8E3512",
            INIT_RAM_11 => X"58AE542A158B05A2FA7D44A351A8DC6860C16CC0A250A34900A30AB75BAED7EB6BCD3469",
            INIT_RAM_12 => X"EB75BCDDEAE73BDDBED6E564702853E9F4EA68B45B4C958A02972279409E312853A5E4C9",
            INIT_RAM_13 => X"8DC6E572B7946E471A853E982F2B2592B7439DC6A251A8542A451A8D42A15128D4AF39A4",
            INIT_RAM_14 => X"B75BAED86BF51564712C964C26130984C2592CA05C5028142A0502813E9F5027D3E9E502",
            INIT_RAM_15 => X"8D48E151A74C09C2E16CAE552904C2E582F27546A472B95C8E04FA95CEE54404D205552B",
            INIT_RAM_16 => X"9148A572295C8E2702D26974BBEE76FB5BC6C6409E4FA8540A04F275369C4E269326651A",
            INIT_RAM_17 => X"8542A05028140A050A95CAE67338140A35228942A04F2AE5B2D9539DC8A65338946A772A",
            INIT_RAM_18 => X"9DD2EC75BADA46874BBB5DAED86C3575E69A34984C26130984B25938B4A371B8D44A3512",
            INIT_RAM_19 => X"793C9E4EA713EA54E974C89D31A85409A30A85409D2883CA2552EA7D46A572B99CAE44A1",
            INIT_RAM_1A => X"A9CEE872A9150E874BA5CEE673B95CAE470A756977DC6EB6B58574A5C8E251A70B861502",
            INIT_RAM_1B => X"5546E673395CAE57238D46A25128146E352B99CAE673399CAE4722853EA04FAA1DD2C95B",
            INIT_RAM_1C => X"8944A573BA1D2E771AA9DB2C97CBA5929743C35FAFD7EC35B658CA449A4D26930984C259",
            INIT_RAM_1D => X"A9C8E14FA68B65B2EA753A9E4EA753CA350A8D3CA053B8D40A050285385D2C164B25A2FA",
            INIT_RAM_1E => X"91429F4FA99E76F96CBA54E874B9DD4EB75CAA4CE874BA1CEE570A60B449090242E69712",
            INIT_RAM_1F => X"591E4D26130964C2818550E873B99CCE672B99C8A573B9DCEE472B9DCEE873B99CCE452B",
            INIT_RAM_20 => X"95385E2C168BC8B2F17D46A673BA9D4EA743B1D2EF97CBE5F2F974C361B0D86C35FAAB14",
            INIT_RAM_21 => X"712E4F070404AE86CA8DB6604EA70C29B2DA813CA04F25CCCE653A8538635227D42A2512",
            INIT_RAM_22 => X"A1D2E674BA5D2E87338540A14F1B26974B74BE5F2E974B656ED96CBA552C954A1CEE050A",
            INIT_RAM_23 => X"BF5FB0D86C35FAED55862A8E26130984C2E2A9D72B74BA5D0E773B99CCE9753A1D0E5743",
            INIT_RAM_24 => X"8942A2522913AA54FA85305F4D160D2DE4A29550E774BA9D6EB753C2673499CCA6733B84",
            INIT_RAM_25 => X"C2DB2E95CA1CAE46F275200E0603050E67437D34604F27D3C9E4FA7D3E9E4FA7540A4532",
            INIT_RAM_26 => X"A1D0EC964AE46CE33BA9D6EB753A9D4E97439546A04F28173B7BBDCAE532984C26132B7C",
            INIT_RAM_27 => X"DEEB76BA5DAE774BA5BB5FAFD7EC35FAFD6DA2BED4471349A5454CBE5D2C963ADD6EB74B",
            INIT_RAM_28 => X"793EA14FA6D3CA655B953C6650A9DC0A151A4CB2614D9921A5A3128546AA753A9D0D34AA",
            INIT_RAM_29 => X"DEE975BADCEE974BBEDF656E954A1CAE050A689E0D0602C50E7712893E9A2F268AE9E4F2",
            INIT_RAM_2A => X"C65F2E96CB65B2C763ADD4EF974A1C2CC34BB2592D964B256EA7439944A150A8973BDDBD",
            INIT_RAM_2B => X"6D1C4A384C25D204C2D6E977BBDDEEF72BBDBB5DAED76BF5FAFD76B2CF1A692389A5C584",
            INIT_RAM_2C => X"893C9D4D971305D4FA793EA05027D38A673A44B29F522A1C4A352299BE9F4F25D205B2C9",
            INIT_RAM_2D => X"9948A25229DDB3ADDEE76B78DCEDF6DB4BB6BA5F6472395C8E24F2549C0D058694EE350A",
            INIT_RAM_2E => X"BB555C6813C9C637A5D2E53098CC2612F973B1D8F197C5D3CCE364B65D2F974B658EB74B",
            INIT_RAM_2F => X"8140A350270C69B2D985C11157CBA651B583E6EF76BB5E2FD9A68ABB5DAED76BB5FAED7E",
            INIT_RAM_30 => X"48220D060B64EE24FA6CBA5D4F268961E4D13C3EA05028142A8732EACAA8743ADCEED74B",
            INIT_RAM_31 => X"C26330984BE5D2D763A9CCA553B8DDF2F9E6D77FFFFCEDF71B6AFBAE4ADE52B95C29E4B1",
            INIT_RAM_32 => X"BB5DAED76BB5FAFD76BB555B6813C9C659B5DAE93299CCE673297CB9E133B8C91CCD155C",
            INIT_RAM_33 => X"A14AA87227946A87433CBE982D178CAA5553A15122774B65D22600C66B78BCDDEF17BDFF",
            INIT_RAM_34 => X"8148DD4B991C2982A9401E0D040A5C6A450A853C9E4EA753A9A2E28140A25128D3EB0922",
            INIT_RAM_35 => X"CA6774B95CECAE499DCEE772B94C65F2E96BB1D4EB712716371B95E36974D75C6FBD834C",
            INIT_RAM_36 => X"206139BEEDEFDF9DE6BB5DAED76BB5DAED76B2CB55489389A669BDDEEF76BB5DAED76BA4",
            INIT_RAM_37 => X"7D3CA25128942A8743B5BA6E869CF54E9722914AD76AAB1C0A053ABE54ED98CD6DB30889",
            INIT_RAM_38 => X"D6EDB1BA5BE429D533693C9E4D96CB0582B94C1E0F0A1B24CE872268BEA14FA81245B2EA",
            INIT_RAM_39 => X"E775BBDD6EB75BADD6DAE967795D6E575BADD6E974BA5CE653097CB9D6E64D960D532BA5",
            INIT_RAM_3A => X"C661319ADCA65192C11406349D6DAF1BBDBEBB5DAED76BB5DAED6EA2B6D0271349A617B5",
            INIT_RAM_3B => X"7D42A150244C09D4F2753C9B31281409C52AA1E928743B1DAE751AADD4DE512914AA755B",
            INIT_RAM_3C => X"C25ADF4E95CBCB4BBECEE32874BA5D0E351A8144982EA70B4592A1502212133A9CEE2512",
            INIT_RAM_3D => X"8E228F269349C57575EB79BDFE6EF75BADCEEB6F72BADD6ED76BBDE2EF76BADD2E933994",
            INIT_RAM_3E => X"A5B0686FA893861573C661329BDCEE3224E2340C001BDEAF9BADE7BB5DADD76BB5DAED6D",
            INIT_RAM_3F => X"64A4121539DD2E66E12C325C2F264BC9D4FA70B45F4E289389D5949558E256BA9D2E0501"
        )
        port map (
            DO => promx9_inst_14_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_13,
            RESET => reset,
            AD => promx9_inst_14_AD_i
        );

    promx9_inst_15: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"DEF3B8BBDDAEB75BACCA50E04FA7936687BED6EB79D8C99C8A350274C0A150A813E9E4EA",
            INIT_RAM_01 => X"B75BADD6EBB5DAFD6D821C4F269349C512F3DB7BFDFEFEF75BCDDEF375B7BA5DEED77BC6",
            INIT_RAM_02 => X"8954E85739DC2AD722CA44A55125DC4A9774CA6777BA5CACAE37026D0E07008DA717ADDE",
            INIT_RAM_03 => X"813EA15028142A04F270BA920F29154E24A114205930A70BCA250275409F4D98938A0502",
            INIT_RAM_04 => X"E773A9954D6EBB4BD6EF75B9DDEE2F177BB5C646A150A813A5B38DEB5D2571A91C8A2502",
            INIT_RAM_05 => X"7D1407040046F79DB5BB5BADD6EBB5DAFD6E7E1E4F269349C502928A6BBDFEFF7F9BCDDE",
            INIT_RAM_06 => X"34286352A38981230ADED2AF78CB1C8A756BA548A55326DC71131CDEEF74BC5CA4EE671B",
            INIT_RAM_07 => X"30C0A15128D429A2F270B65D4F26CBE9E4FA7D3E9E4C9A5D4E76A2512E5F50250BE86102",
            INIT_RAM_08 => X"4D40F1BDEF7F9BADADBED12ABBEEB6DB9DF7F7FBFCDDEEB75B8BBDA9C8A15127D3E9D2E1",
            INIT_RAM_09 => X"E773B7BAD99D0E7723853686040200A39BBDBF5DAED76BB5FAFD6E92248F271349C4F289",
            INIT_RAM_0A => X"24B05E53330C8D04594022582D124164B2FA70D6F09D5C64EB0722A9D2A14F27DBEEEBC5",
            INIT_RAM_0B => X"914CA551A813E9E4EA28BCA052381409E4D960B49D4B95CBA5C4E18942A14E1ADDD296D2",
            INIT_RAM_0C => X"A2B291279349A4E27944A69B5249E4B226EB652A9B744A65938DCEE375B8DE6EF77BAD84",
            INIT_RAM_0D => X"9D58EB92CAEE97ADC6EF6D6F8F2AE52E97338DBA8904824140C240BF5FAFD76BB5DAFD6E",
            INIT_RAM_0E => X"7142A350AC6653184024C6A76996D261F4F28146A351299C6C80CA9DBCBFDA4D264F0742",
            INIT_RAM_0F => X"D6E52F963ADD2E87329D4EE652289429D2A254C0A14F264B69C4E2752C582D944A04C068",
            INIT_RAM_10 => X"BB5FAFD7EBB5DADD6EAAC313489389C4D2713CA2522924D2A954AA55289229144ACAE9B5",
            INIT_RAM_11 => X"554ADE5FFA1717ADB4E6E734B95E377B6BD6C2D72A954B250E87338DBC8D04024140B061",
            INIT_RAM_12 => X"68B6480D94CB89E4E28544A3502C6E5185AE28B4634916CCCE452A7940A15129DD0E4669",
            INIT_RAM_13 => X"44A250279389E627BDDEE97096BB5D6E9743A9D0E77329142A96EA853A9B2FA64A65A2D9",
            INIT_RAM_14 => X"8DBC8904028140B061BB5DAFD76BF5DADD76AECF5E6B24D204E271349C5028948A453492",
            INIT_RAM_15 => X"9DBCA25439DC4902916D4ECE2AAC6FDF8BD5F373B7BDEDEEFB6DB5B65B2D964AE552A93B",
            INIT_RAM_16 => X"7124192D16CB85A2B950AE5A2E150BC9F50A7D42A153BDE86196AA34AC9E532A5CCE7743",
            INIT_RAM_17 => X"409E4E2793CA04F2793C9E4F271389C5658DE6ED7196BADD2E9753ADD8EA7439948A14FA",
            INIT_RAM_18 => X"BA34AD97CC2DB2B9448DBA8704828164C261BB5BAED76BB5FAED7EB75768B1C79B6D749A",
            INIT_RAM_19 => X"552AA151A7D50E974BA1B46453BA9D5204FAA1D2C90692CD8E974BB6571E56DCEE76E984",
            INIT_RAM_1A => X"B1DF2F96CA1D2E670A60A65A2D154AE582A960B2582B174BA9F4E18148A7722D6AA9F6DB",
            INIT_RAM_1B => X"BF5DABB55AAD768AE34D1E4E271389C4E271389C4D269389C4F31BE2F173B84B654E4743",
            INIT_RAM_1C => X"DEDF33B9DC6D56E9239650F0B7CBA5B2B93385B48804828160C261B35BADD76BB5FAFD7E",
            INIT_RAM_1D => X"852C4D1026CE1248AA9DA269753A9D0E874BA1D8EC7537114686DAAE54E24592CD52E964",
            INIT_RAM_1E => X"C2F174B7C85C0ED953AE653398CADDB2871A5CA6592903C20100784C2E5C2E191161E4F2",
            INIT_RAM_1F => X"AAD76CB66B75DAFD86C35FAED65B2D96CB1449204E269389C4E271389C4E271349C4D2BA",
            INIT_RAM_20 => X"AE54DA4613CB2AF96589DB2F99DBAD55555469A4AB96CB65F668BA6D224804828184C269",
            INIT_RAM_21 => X"5CB04C2688544992FA8536624603C716997CCE5CEA763ADDCEB753A1D4E656CB279EC90B",
            INIT_RAM_22 => X"349A4E269389A4D27181EF79D4469CD3296CB66532974B1BCA971A5CAA6468971B256280",
            INIT_RAM_23 => X"288E0704828184B261A6D56BB5DB2D96ED7EC35FAFD6EB2DB6CB1C4D1E4E269349A4D269",
            INIT_RAM_24 => X"ADD4EC9B6CAD92CAC3AE571344034C730BBD7E4EF4B9DE34B4F52524D52C95CB253256AA",
            INIT_RAM_25 => X"9DC29844186325111B5CB25E4E970BA9D5128D36624E181306579DD2D8EE774C2632B75B",
            INIT_RAM_26 => X"449E4D269349A4D269389C4D269389A4D26940CF37B54AA6972954A9DF3197CADC2E1522",
            INIT_RAM_27 => X"C6BCE893CAE4ACE282248E090502C964C2619AD169B55AAD76CB6EBF61B0D7EBB5BADB1C",
            INIT_RAM_28 => X"6958EC784A5C0D455B99F1B1964B6573097CB6592165999EBBFFAEFBC527774CEE5BFFFF",
            INIT_RAM_29 => X"CEE32C97499E571953ADD8E56A250A05035CBA345A2D9893EA54EA81366150A344CF3995",
            INIT_RAM_2A => X"BB5FB0D86BF5DADD1C409C4D269349A4D269349A4D271349A4D26934AAAA9CEDEF174B94",
            INIT_RAM_2B => X"DF77FDF85DB6562734A2472072395C0D126120100904824184C26996CD67B45A6D56AB66",
            INIT_RAM_2C => X"70C8A152A9558E15CDC2613399DD2A89657CB65D30B8DDEE379D94BA5D2D86934E772B95",
            INIT_RAM_2D => X"349C57554E773B5BBDDAED667849E42F198CBE54E970AA9D2EA72BDAB66250AA1C2A5533",
            INIT_RAM_2E => X"96CD67B3DA2D169B5DB6DDAFD7EBF5FAED24409C4D269389C4D269349A4D271349C4D269",
            INIT_RAM_2F => X"C261309BE9A6178DDED2DF2EB8DBA79F8F34CADD2B94485A65023820120A0502C984C269",
            INIT_RAM_30 => X"C65D2671299C8A6753B1CEEE99CCE612D9D6E76535BD6B22EB28AACADF31BA5CAEB70B8D",
            INIT_RAM_31 => X"349A4D269349A4D269389C4E2AAA671B8DC6E36F6B995CAE9B7B94CA52EF96B8552F2953",
            INIT_RAM_32 => X"20140B2502C984C26996CD67B45A2D168B4DAED96DD76BB5DAED34449C4E271389C4D271",
            INIT_RAM_33 => X"CAED73BADD6E574B8DCAE139D4CE76DB5BC6BEF7F7DD728F7B0B9DBA5925713712A48048",
            INIT_RAM_34 => X"D6DF30994A9CAAE9B5BA54E773B8D4AEC712BE676C953DEE96E96CF36576BA571D519459",
            INIT_RAM_35 => X"491C4E271389C4E269349A4D269349A4D269389A4D26944C4F4BDEEB7177DB6E767659CD",
            INIT_RAM_36 => X"B255206D250920904824144C25930984C27996CD67B45A6D368B45AAD76DB6EB6DB6DB3D",
            INIT_RAM_37 => X"EF3AF6BE6208E156A2CAFBEF9C6DF6FB4BA5D2EB647039A79F5D24DB6B73BF7FFCF2D97C",
            INIT_RAM_38 => X"EB77B8DBEDF71ADBA5DEEF7499CCA633AB94C6306C753A9D0F196CB6632477C89EB72984",
            INIT_RAM_39 => X"A6D56CB6DB75BADB354D1E4E271389C4E271349A4D269349A4D269389A4E271389C59554",
            INIT_RAM_3A => X"F3FBEDB8DCAE570B0B99BC9326924120A0502C964C269309C4F27996CD66B3DA2D168B45",
            INIT_RAM_3B => X"C66575BADD2F9B2B84C6556EBCE5128924BBDF73B6DDEDF6FBBDADCECAE56B2D35976DD7",
            INIT_RAM_3C => X"349A4D269349A4E2817DE37BDE7EB71B5D75DEEF76B9CF36B75B8CD2CEF192AB1D2E97A4",
            INIT_RAM_3D => X"9ECF66B359ECF67B3DA2D36BB6DB6DBADB4D5D1E4E271389C4E271389A4D269349A4D269",
            INIT_RAM_3E => X"95D0E673385EDBBFD7B2576B99DAA532670361264905028140A051309A4D271389E4F281",
            INIT_RAM_3F => X"E6CF39B84C65B3096BCA6D78BADD2E974BC5BA267FFB5D75136D2CDB7BFBDEFF7EFB7D9D"
        )
        port map (
            DO => promx9_inst_15_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_15,
            RESET => reset,
            AD => promx9_inst_15_AD_i
        );

    promx9_inst_16: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"83C1D8CC6633198A8562B198CC6433198CC563026B8A692D99CCA5D037C9D142855AB014",
            INIT_RAM_01 => X"2131188C582C160B4696BAD5469349A4D269352AE596ED7FBFE16C6CC1E110883B1D8EC7",
            INIT_RAM_02 => X"8EEB433A3EF05EAE4824F27974A03D100083419171C4AA2A1203C0E0F0783C2E08088643",
            INIT_RAM_03 => X"2E4713B2C55C592BA4708783F56DAD6428D6ECE5AAD15AAE5EB5D224815156235A6824DB",
            INIT_RAM_04 => X"50626110763B1D8F078431D8EC6633198CC662B198CC6633198C85633160BD00FC83C5A1",
            INIT_RAM_05 => X"E08080202211108683623158B05834168D46D7DB9D8AA349A4D269352A954AB964B6DCEC",
            INIT_RAM_06 => X"4022F0A464FA982ED88E966B156CB2768D0FA792C098B43D130300A06070180E0F0785C1",
            INIT_RAM_07 => X"62B198A8562D1A1B0D4402045E60FDC55BB23249DDF661196FBB4EAA754B017CB86F35CA",
            INIT_RAM_08 => X"34FA0506934AA954AAF354E910783C218EC763B1D8EC783C198CC6633158CC6633198CC6",
            INIT_RAM_09 => X"A050383C101004020101108844241B1106C4624160B05A2C168D46197C2DF2C559A8D469",
            INIT_RAM_0A => X"2686BC21A6E369A315075000B890052506CCE262826CC8723690CE4682F9349A23060300",
            INIT_RAM_0B => X"633158CC5633158C85632190A8542A150AC462C160A4854197C7D736D73315D4038D3ED7",
            INIT_RAM_0C => X"5A1C863AFB74B1D66A348A34DE7F3FA0D2AA3498315488441D8EC763B1E0EC763B1D8CC6",
            INIT_RAM_0D => X"E87159C46A19060100A070405C101008044321A0D06C462411890582C170D46A2D1A8D46",
            INIT_RAM_0E => X"D1D6A6562A00AC39574F3872A85C1500218D8844B9EDC9C950A98DE7746C8DD02C5A1600",
            INIT_RAM_0F => X"63B1E0F0783B1E0EC6833190AC6633158C8542A150A8542A150A8542A150A854203D376C",
            INIT_RAM_10 => X"C361F0D87A361F0F87BB3D5EAB3197C2DD2D559A85228F3FA050AB557982DCA8441D8EC6",
            INIT_RAM_11 => X"423562C104A45F238F02233960781B068180E1004040201108864241A0D09058251A0B45",
            INIT_RAM_12 => X"42A14888542A1088D6D19933E9CA9A3F2A0FACD1E91C240000B760492358481972331C0D",
            INIT_RAM_13 => X"347A142CFC55218EC642A198CC78451E0F06633198CC562B198CC542A158A8542A150AC6",
            INIT_RAM_14 => X"6221106C461E1F0D87C361B0D46C361F0F87FCEE2EF779AAD0E431D7DB9D8EB551A45028",
            INIT_RAM_15 => X"4DF2A2E0A69233FEA08B760A4952514B21906712D93048060383C1008040202210088483",
            INIT_RAM_16 => X"42A150A8542A150A8542A150884222108845F0CA4CFA68B68020CD04C1C8A80A0202BE19",
            INIT_RAM_17 => X"398C861EFB6BACD429147A2CB5B4762A90C7432150CC663B1E1107834198AC5633198CC5",
            INIT_RAM_18 => X"0110884434220C848362311890482C168D87C361B0D45C3E1B8F861D7E7F3B8DC5DE6CF5",
            INIT_RAM_19 => X"42E088181C0D02BA5B4DD1BA6A50EA7BF7EC5AF6B1E994EA4C2191475278B40E06038201",
            INIT_RAM_1A => X"83C1E0CC6633158CC642A150AC542A158A8542A1508844221488444272ACC5809F4410C6",
            INIT_RAM_1B => X"FC8EBF3F9FCFE36F779B3D5E87218EBADAAA349A44F238D13712C7632150C86432198D07",
            INIT_RAM_1C => X"E621381C0E080402012120C848341B1106C462311890582C120905C351B0D86A361B0D86",
            INIT_RAM_1D => X"22110054423A1C8803A16028181A070700DD4A9683762F49C7C5F7E5879AC1EAC3569F90",
            INIT_RAM_1E => X"83B1D8C8542A150A866331D8CC6432190C8542A158CC6632150A854221488854290C8844",
            INIT_RAM_1F => X"823128B05A2D1B0F87DCFE7F3F8FC7E36FB7DBDDA6B35599CBE1AEB6BAD542891C699F8A",
            INIT_RAM_20 => X"DAFE7DBD008F47224CA0803800100804824241209068361B11890582C1208C4623120905",
            INIT_RAM_21 => X"422110A8542A1488442211088040180F85C2E17070380E0F0405808FE5D3B6E35AC270F5",
            INIT_RAM_22 => X"F7DBA5AEC5579CBF1005D258E86429148A8542A158C8542A150A8442B160D06632150A85",
            INIT_RAM_23 => X"62412090582C16090582C160B0482C158B059B5DEF1B8DBEDF6FB7DBEDF6F769ABD0E431",
            INIT_RAM_24 => X"00F60349F7138DCC708EE733BD8E864AA00000804020120904848341A1186C361C1186C4",
            INIT_RAM_25 => X"42B1A0CC642A150A8542A150A8542A11088542110860301F0B85C20180B8202E08080242",
            INIT_RAM_26 => X"BBEDB6FB7BB4D5E8B238FC3DFAEB6BB0D3224B33F1508633190A85429150A45221108A85",
            INIT_RAM_27 => X"61B0D88C482C1208C462312090482C160B0582C1208C4623120AC55ABD9ED37BBEDF6F77",
            INIT_RAM_28 => X"0180886420110C0402010098AA13418B4EA4930AD3B1749530824120908024120A090484",
            INIT_RAM_29 => X"432150A45229150AC6633198C8542A150AC662A150A8542A150A842211088440180C0602",
            INIT_RAM_2A => X"39AD5EAF59B4DA6D769B5DAEDB6DBEDEED34799C461EFD75BADD2C34283A8CF05E2610C7",
            INIT_RAM_2B => X"4120904C3412090483624120AC4824160904824120B05824160B0582C1608C482B120B05",
            INIT_RAM_2C => X"2211088442180C86030191088430110C04020110904C424887381E1535F2F97612050281",
            INIT_RAM_2D => X"D73ABCD6491874AA8EE572B1349C572F1548A42148A85633158CC642B158C8542A150A44",
            INIT_RAM_2E => X"82C160B0582B158AC5191CCE8B45A3D66B359B4D6ED35BB5DB6F759AACC63EFD7EBBDFEF",
            INIT_RAM_2F => X"67A3984C26130984826130D86C361B0D88C4824160B0582C160905624158B0582C160D05",
            INIT_RAM_30 => X"42B198C8542A14888442A1108442211088442211088444211084422190E0A83A230D058C",
            INIT_RAM_31 => X"9ABD0E230187BFE030187BA56EB963B15469F3591C45F0F1792E8EE4A148A8562B198CC6",
            INIT_RAM_32 => X"62311088382C160B05A34160B0582B158AC5190C8E67339AD168F59ABD5EB359ADDAED76",
            INIT_RAM_33 => X"21B150AC4A2C1188C461B0D86C361C0D86C261B09870482411870582C168B45A2D168B05",
            INIT_RAM_34 => X"05B190AC6633198CC6633198AC662A150A8542A150A85421108844221100644221110844",
            INIT_RAM_35 => X"39AD168B47A4D66975BB4D16471388C4E231185BA592CB6EBF5FAEB74B65B2DB74B1559C",
            INIT_RAM_36 => X"82C168D46A351A8B46A320E0AC441D198905834160B04623160D05190C8E673399CCE673",
            INIT_RAM_37 => X"2211088442200C8844221110B05C35120AC461C12090381C0E06C3824128B04824128B05",
            INIT_RAM_38 => X"B75BADDAFD7FC2DBE8063198AC6633198CC6633198CC6632150A8542A150A85422108844",
            INIT_RAM_39 => X"198C86633398C86432190C8E67359ACDE7359ACD5E8F359AC8E27118FBEDB2CB76BF5DAE",
            INIT_RAM_3A => X"A2D160945824128B05825168B45A2E1A8B05A2C128D46624160B0582C160B4582B160CC5",
            INIT_RAM_3B => X"62B150A8542A150A85421110844221108844222150B06C35160945A2D160904A2E1A8B86",
            INIT_RAM_3C => X"187BEDB6EF87C3E1F0D7EBF5FAEB75BEDEAB684198AC6633198CC662B198CC5633198AC5",
            INIT_RAM_3D => X"82C160B0582C1A0B05198CC6432198C86432F90C8E673399CD66F49ACD66AF459AC8E471",
            INIT_RAM_3E => X"A2D168B04825168B8604E1B0D46C35168B868220E8B45A2D1A8D4682D168D4682C1A0B05",
            INIT_RAM_3F => X"633198A8562B198A8562B150A85422150844422150844221108885222150B06C35168B45"
        )
        port map (
            DO => promx9_inst_16_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_17,
            RESET => reset,
            AD => promx9_inst_16_AD_i
        );

    promx9_inst_17: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"389C4D269349A4D261349A4D269349C4E27138A6A89AEE371B7DAECAF5B5BCDCEEF76BA5",
            INIT_RAM_01 => X"309C4E2713C9E50289A6D167B359ACD66B359ED169B55B2DB6DB556D9C4F271389C4E271",
            INIT_RAM_02 => X"E77DF6DDEDEEDB4B4CAA50E772381BA9027138AAA36FB6D309225824140A05028164C261",
            INIT_RAM_03 => X"BAE379DEFF3EF74BDEE773B9D6CFBED71BA5E6F176BADD6ED75B8475D71D7F6C75F6ABCE",
            INIT_RAM_04 => X"86204E271389C4E271389C4E269349A4D269349A4E269349C4D269389A4E2D2AAE174B95",
            INIT_RAM_05 => X"28164B25930984C269389E4F27940A050289AAD569B3D9ACD66B359ECF67B45A6D56BB4D",
            INIT_RAM_06 => X"30D71C54CEB7DF6DCEEB6FB4BA5D2EF96564B6532072B81B8952381C120904828140A050",
            INIT_RAM_07 => X"389C4E26938A0564BA552AB4DDEDB7DFEFFFDF75BDFDEE76BB7B84DAF178DB6D2EFB4B43",
            INIT_RAM_08 => X"9ACB25B359ACF68B4D962E8F271389C4E271389C4E271389C4D269349A4D269349A4D271",
            INIT_RAM_09 => X"20100A0502C964B2592C984C261349A4C2713CA04F27940A051289B3576AB4DA2CF67B35",
            INIT_RAM_0A => X"AE73BCDB6E76575BB57A0E196F34938D44DB613CEEB4CB25522754AA5325723712651238",
            INIT_RAM_0B => X"349A4D269349A4D269349A4D269349A4D269389E4F2AAFFE5AFB6CEFE975B955173B6DA5",
            INIT_RAM_0C => X"BB5BACD5DAAD568B3D9ACB6492C964B27B459AC111279389C4D269389C4E271389A4D269",
            INIT_RAM_0D => X"BA2AAA90375328804020140B2502C964B261309A4D271389C4F28140A05128940A251289",
            INIT_RAM_0E => X"EB6974D5D2CFDF5DA5E775AE8DA5C9E33B8C8A411D74DEFC7208E3B65F3BD556DE557672",
            INIT_RAM_0F => X"349C4E271389C4E269389A4C269349A4D269349A4D269349A4D269349A4C26134B6EFBF7",
            INIT_RAM_10 => X"40A25129144A451289C75FAFD76B7596BB4DA2CF66B2D964B26B45A2C91A6893C9C4D269",
            INIT_RAM_11 => X"79E573B75C2E76D96475D1267036D100905028164B2592C984C261349A4D2793CA04F279",
            INIT_RAM_12 => X"30984B26130984B344CEEBB2B458A512F954B63E9E4C94C8C39DDEAABF1048AFBD11D6EC",
            INIT_RAM_13 => X"9ACB218AA409C4D26930984D271389E4E271349A4D269349A4D26930984D26130984C269",
            INIT_RAM_14 => X"349C4E27938A25028940A05128944A451289CF67B1D8EC35FADD66AAD569B459ECF66B2D",
            INIT_RAM_15 => X"EB3AEAAF4CEBCFFFB6CAED70B85A2616E96CAA51226DA20120A0582C964B25930964C261",
            INIT_RAM_16 => X"30984C26130984C26130984C2612C984B261AA6DB5D7D9A676991B85B89A4A1300C3CDB6",
            INIT_RAM_17 => X"BB5BADD65AAD167B359ACB248EB55224F26930984C269349A4E271389C4D269349A4D269",
            INIT_RAM_18 => X"2C984C261349A4C269389E4F2793CA05028944A25027948A252289D7E7B3D9ECB65B1D7E",
            INIT_RAM_19 => X"6D2E52260241433BBEE33CE59EFDF6FBFFD6EFEB6E97DE3616FB74AA48DE44828140B059",
            INIT_RAM_1A => X"389C4E269349A4D26930984C26930984D26130984C26130984B25930A26FB24964ADF6DA",
            INIT_RAM_1B => X"D369F4DA6CF67B2D96C761AFD76B7596AB459ECD65B1C75AA9027134984C26130984D271",
            INIT_RAM_1C => X"99B08905028164B26130984C269349A4D271349E4F2793C9E4F28140A05028140A251289",
            INIT_RAM_1D => X"2C964A2815530984B24C960904824140A1C6C6EFB6DC6E375F0BF785EBB3BB6CEE36B964",
            INIT_RAM_1E => X"389A4C2612C964B261309A4D26930984C26130984D26934984C26130984B26130964B259",
            INIT_RAM_1F => X"3C9E502813CA251289CF69B3D9ECF67B2D96CB65B1D86C35DADB5DAAD367B35923AD5489",
            INIT_RAM_20 => X"F7FBFAD74BADD2D95448964B05930984C269309A4D269349C4E271389E4F2793C9E4F281",
            INIT_RAM_21 => X"30984C26130984B2592C964B25128944904828120A04828140A250E76976DFFF3F7FDFE7",
            INIT_RAM_22 => X"B2D76AB4DA6CD228B2491E4D26130964B25930984D26130984C261309A4E27134984C261",
            INIT_RAM_23 => X"389C4F2793CA04F28140A04F2793CA04F281C363B2D96CB65B2D96CB67B2D96C761AFD76",
            INIT_RAM_24 => X"30D535DB6DB6BB6DD7BEE374BADB65B2B869309A4B261309A4D271349C4E269389C4D271",
            INIT_RAM_25 => X"309A4E26930984C26130984C26130984C26130964B25128920904828944A05928164B259",
            INIT_RAM_26 => X"CB65B2D9ECB65B1D7EBB5B6DB5DAAD369B2471AA9127934984C2592C964B2592C964B261",
            INIT_RAM_27 => X"389C4E2713C9C4F271349C4F2793C9E502813C9E4F2793C9E4F279BB5FB0D8EC765B2D96",
            INIT_RAM_28 => X"28944B2592C984B2592C984F3AEF3E9B9DAEDF73F6D9DC2C4CC269309A4C261349A4D271",
            INIT_RAM_29 => X"34984C2592C964C269349A4D26130984C26934984C26130984C2612C964B25928944A251",
            INIT_RAM_2A => X"B35DAFD7EC363B1D8EC763B2D9ECF67B2D8EC35DADD65AED76BB5DA6C71A4B245204E269",
            INIT_RAM_2B => X"389A4D271349A4D271389E4F2713C9E4E271389C4E2793CA05028140A04F2793C9E4F279",
            INIT_RAM_2C => X"2C964B2592C944B25128964B2612C984B2592C984D2795167B1B9EEBDF71BA5409A4D269",
            INIT_RAM_2D => X"B6D56793496431A6AA44A05028140A2502793C984B261349A4D269309A4D26130984C259",
            INIT_RAM_2E => X"40A050279409E4F279B359ADD76BB5FB0D86C763B1D96CF67B3D9ECB61AED6DB2D96DB6D",
            INIT_RAM_2F => X"7DBACE271389E4E269389C4E2713C9C4F279389E4F2793C9E4F279349C4E2713C9E50281",
            INIT_RAM_30 => X"309A4D26130984B26130984C2592C964B2592C964C261349A4D26130984F269409E4E2CA",
            INIT_RAM_31 => X"CB63AED6EB75B6DB76B7596AB4DAAD569B4D9E4B249148A471B6AA44984B261349A4D269",
            INIT_RAM_32 => X"38984D269389E4F279409E502813C9E4F279B359ACD66B75DAED7EC35FB0D8ECB65B3D9E",
            INIT_RAM_33 => X"309C4D27140A04F279389E4F2793C9E4E2713C9C4F2793C9E4E2793C9E4F27940A04F279",
            INIT_RAM_34 => X"491A4C269349A4D269349A4D26934984C26130984C26130964B2592C984B25930984C261",
            INIT_RAM_35 => X"BB5DAFD7EC363B1D96CF63AFD7EBB5DAED76B7576AB4DAAD76CB5DAED56BB5DB2D768AF3",
            INIT_RAM_36 => X"3C9E5027940A05028140984E269309E4E27940A0502793C9E50281B359ACD6EB75BAED6E",
            INIT_RAM_37 => X"2C964B26130964C25930984D27944A0502793C9E4F2793C9E4F2793CA0502793C9E4F279",
            INIT_RAM_38 => X"AAD56AB5DB2D96AB2C4D1C4D269349A4D269349A4D26934984C26130984C26130984B259",
            INIT_RAM_39 => X"B359ACD66B359ACD66B35BADD76BB5FB0D96CB65B0D86C35FAED76BB596AB4DAED76BB55",
            INIT_RAM_3A => X"40A04F2793C9E4F2793CA05028140A0502793C9E4F279389E4F279389E502813C9E50279",
            INIT_RAM_3B => X"349A4C26130984C26130984C26130964B26130984D27944A25028140A04F27940A24F281",
            INIT_RAM_3C => X"BB596AB5DB2D96CB65AED76AB55AAD56AB45511A4D269349A4D269349A4D269349A4D269",
            INIT_RAM_3D => X"389E4F28140A04F279B359ABD5EB759ABD66B2D9ADD6EBB5DAFD86C765B2D86C35FAFD7E",
            INIT_RAM_3E => X"44A25027940A0502894D225128140A0502813C9A5027940A0502813CA04F2793C9E4F279",
            INIT_RAM_3F => X"349A4D261349A4D261349A4C26130984C25930984B2612C964B261309A4D27948A251289"
        )
        port map (
            DO => promx9_inst_17_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_17,
            RESET => reset,
            AD => promx9_inst_17_AD_i
        );

    promx9_inst_18: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 18,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"B6FC2BBF0AEFBEBBF0AADBEAB6EA6CBA7AAB65958E30734B18D2C634B18D2C634B18D2C6",
            INIT_RAM_01 => X"C74D32D35C74D70CF3BF2CEFCB2BB1C6DC31B6FC2BBAEAACB2AB6DB2FBECBF0B2FC2CBF0",
            INIT_RAM_02 => X"B30CEBBF2AEFCABC32AF0CABBF1AF0CACC32B30CADC33B70CEDC73B71CEDC72BB1CF0CF4",
            INIT_RAM_03 => X"40D18F3053CD18F34638B10F3463CC14F3053CD14E3053CC14F3053CB14F3053CC150305",
            INIT_RAM_04 => X"40D19034644E19038640D19034544E19034644E18E2C440D14F34540D19034640D190345",
            INIT_RAM_05 => X"30A14D28534B18E30544E19138644E15138644D15134544E15034540D15034540D150346",
            INIT_RAM_06 => X"30A14D2C530A14D2C530A14C28530A14C28530A14C28530A14A2032880CB2442C910C284",
            INIT_RAM_07 => X"71D70F34834B18D2C634B14D2C634A18D2C630A18C28534B14D2C630A14D2C534B14C285",
            INIT_RAM_08 => X"B2FBEAB6DA2BAE9B2CAEEBABBF0AEFC2BBAFAAEBEBBAFAEFBEBBAFAAEBE9B2EA2CBA7AAC",
            INIT_RAM_09 => X"B70CADC32B70CEECB4BB2D2ECB3BB1CEFC72C33D31CF4C33D30CB4BF1CEFCB3BB0C6DC31",
            INIT_RAM_0A => X"3CD18E30538C10F3053CC14F3463CC14E305B30CECC33AEFCABBF1AAFC6ABB1AEFCABC32",
            INIT_RAM_0B => X"44E19138644E18E30440D1503463CD15038640D19034540D19034640D18E3043CD14E305",
            INIT_RAM_0C => X"40D15138544D19138544E19138644E19138644E19038640D19034640D19038640D150346",
            INIT_RAM_0D => X"30A10C28530A14B2442C910C28430A14C28430A14D2C634B14D2C634C14F34638B14E305",
            INIT_RAM_0E => X"34B1CD2C634B14D2C634B18C28530A14C28530A14D2C530A14D2C630A14C28530A14C285",
            INIT_RAM_0F => X"AEEBEAB6EAADBEAB6FAAEC2AB6FA6CBA8B2D8638D138934B1CC28630A18D28634A18D286",
            INIT_RAM_10 => X"BF1CB0CF4C32CEFC72BF1CAFC72BF2CAFC72BB0C2BB6DA6BB29AECAADB6BBAFAEEBECBAF",
            INIT_RAM_11 => X"B30CECC33AF0CABBF2AAFC6ABB0AEFC6BBF2AEFC6DC32B30CADC72B71CADC32BB1CEDC72",
            INIT_RAM_12 => X"40D19034640E1903463CC14E2C43CC14F3453CD18F30538C14E3043CC14F30538C14E2C4",
            INIT_RAM_13 => X"44E19138644E1D138744E1D034640D15034640E19034640D19034540D19034640D190346",
            INIT_RAM_14 => X"30A14D2C634B18D2C634B18B24430A14D2C634A15034644E19138544D15138644E191386",
            INIT_RAM_15 => X"30A14D2C530A14D2C534B14D2C630A14C28530A14C2852C90CB2442880CB2442C910C285",
            INIT_RAM_16 => X"9A9A5340B3CD20D2C634A18C28634A18D2C734A18D2C734B1CC28634B18D2C634B18C286",
            INIT_RAM_17 => X"BF1C6DBEFAACB6AB6DAADBABBAFAEEBEBB6EAEEBEAB6EA6DBE9B6EAADBEABAFAADBE9B6E",
            INIT_RAM_18 => X"AEFC6CBF1AEFC6CBF1B71CADC32B70CADC72BB1CAFCB3BF2CEFCB3BB1CAFC72C32CB0CB2",
            INIT_RAM_19 => X"3CD18F3453CC14F3053CC14E2C438B10D2C4AF0CEBC33AF0CEBBF2AEFCAABB1AAFC6BBF2",
            INIT_RAM_1A => X"40E19034540D15034640E19034640D1903463CD15034640D15034640D18F34630A0CF346",
            INIT_RAM_1B => X"34B18F34644E19238640D15138648F1D238648E19138644E1D034640E19038644E1D1386",
            INIT_RAM_1C => X"30A10C2842C910B24528810C24430A14C28530A10C28534B18C28530A14C28530A14E307",
            INIT_RAM_1D => X"34A18D28634A18D28634B18C28630A18C28630A14C28530A14C28530A14C28530A14C285",
            INIT_RAM_1E => X"AADBAAB6EA6DBA9B6FAAEBEAB6FAADBE9B2F9AAAD861540E24D2C734A18C28630A18D286",
            INIT_RAM_1F => X"BB1CAFC72BF1CAEC72BB0C6EC71C32CF0CF3BF1CADBF0AEDBABB6DB2FBEBBAFAEEBEBB6F",
            INIT_RAM_20 => X"AAEC6ABF2AEFCABBF2AAFCAABF2AEEC6BBF2B30CACBF2AEEC6ABB0AEFC6CC32B70CAEC72",
            INIT_RAM_21 => X"40D1503453CD1503873CD1903463CD18D2C338C14D2C43CC14F30538C14E2C438B10E2C4",
            INIT_RAM_22 => X"48E19138648F1D23C844E19038644E19038644E19138640D19034540D19034640E190346",
            INIT_RAM_23 => X"34B18C28534B14C28530A14C28434B18E30734B18E30648E19134544E19238644E191386",
            INIT_RAM_24 => X"34A18C28630A14C28530A14C28530A14C28530A10B2852C914B2442C910B24330A14C284",
            INIT_RAM_25 => X"9EBB5F86140E24D2C734A18D2C634B18D28634B18C28634B18D2C634A18C28634B18D286",
            INIT_RAM_26 => X"BF1C6CBAFAEDB6BBAEB6FC2DC30B6FC2CBEFAADBA9B2EA6DBE8B2EAADBEAB6FA6CBA9B6F",
            INIT_RAM_27 => X"AEFC6BBF1AEEC6ABB0AEEC2CC31B70CADC71B71CAEC72BB1CAEC71BB1C6EC31BF1CB0CB2",
            INIT_RAM_28 => X"3CC18C28334C14E2C534B10C24238B10F3059ECBE9B70A6EC6ABF2AEFCAABF2AEFCABBF2",
            INIT_RAM_29 => X"44E1D138644E1D034544E19138640D19038640D1503463CC15034540D18F3463CD150387",
            INIT_RAM_2A => X"38C18E30640E19138648E19238644E19138644E1913864CF1D038648F21138644E190346",
            INIT_RAM_2B => X"2C914C2452C910B2042C910B2442C910D2C530A14C28530A14D2C630A14D2C638C1CE306",
            INIT_RAM_2C => X"30A18D2C734B18D2C634A18D28630A18C28630A18C28530A14C28434B14C28530A14C285",
            INIT_RAM_2D => X"B2FC2AB6FAADBE9B2FA6CBA9B2EAADBE9AEEA2BBA49E940D28F34934B1CC28630A18C286",
            INIT_RAM_2E => X"BB1C6DC31BB0C6EC72BB1C6EC71BF2CAFCB2BF1C6DBEFAEEB6CBAEB70C2DC31B70C2CC30",
            INIT_RAM_2F => X"9EBBA7B2FA2CBE9B70AAEC6ABB1AAEC6ABB1AAEC6ABF1AEEC2AB6FAAEC2BBF1B70C6DC31"
        )
        port map (
            DO => promx9_inst_18_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_19,
            RESET => reset,
            AD => promx9_inst_18_AD_i
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ad(14),
            CLK => clk,
            CE => ce
        );

    dff_inst_1: DFFE
        port map (
            Q => dff_q_1,
            D => ad(13),
            CLK => clk,
            CE => ce
        );

    dff_inst_2: DFFE
        port map (
            Q => dff_q_2,
            D => ad(12),
            CLK => clk,
            CE => ce
        );

    dff_inst_3: DFFE
        port map (
            Q => dff_q_3,
            D => ad(11),
            CLK => clk,
            CE => ce
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => promx9_inst_0_dout(0),
            I1 => promx9_inst_1_dout(0),
            S0 => dff_q_3
        );

    mux_inst_11: MUX2
        port map (
            O => mux_o_11,
            I0 => promx9_inst_2_dout(0),
            I1 => promx9_inst_3_dout(0),
            S0 => dff_q_3
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => promx9_inst_4_dout(0),
            I1 => promx9_inst_5_dout(0),
            S0 => dff_q_3
        );

    mux_inst_13: MUX2
        port map (
            O => mux_o_13,
            I0 => promx9_inst_6_dout(0),
            I1 => promx9_inst_7_dout(0),
            S0 => dff_q_3
        );

    mux_inst_14: MUX2
        port map (
            O => mux_o_14,
            I0 => promx9_inst_16_dout(0),
            I1 => promx9_inst_18_dout(0),
            S0 => dff_q_3
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => mux_o_10,
            I1 => mux_o_11,
            S0 => dff_q_2
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => mux_o_12,
            I1 => mux_o_13,
            S0 => dff_q_2
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => mux_o_15,
            I1 => mux_o_16,
            S0 => dff_q_1
        );

    mux_inst_20: MUX2
        port map (
            O => dout(0),
            I0 => mux_o_18,
            I1 => mux_o_14,
            S0 => dff_q_0
        );

    mux_inst_31: MUX2
        port map (
            O => mux_o_31,
            I0 => promx9_inst_0_dout(1),
            I1 => promx9_inst_1_dout(1),
            S0 => dff_q_3
        );

    mux_inst_32: MUX2
        port map (
            O => mux_o_32,
            I0 => promx9_inst_2_dout(1),
            I1 => promx9_inst_3_dout(1),
            S0 => dff_q_3
        );

    mux_inst_33: MUX2
        port map (
            O => mux_o_33,
            I0 => promx9_inst_4_dout(1),
            I1 => promx9_inst_5_dout(1),
            S0 => dff_q_3
        );

    mux_inst_34: MUX2
        port map (
            O => mux_o_34,
            I0 => promx9_inst_6_dout(1),
            I1 => promx9_inst_7_dout(1),
            S0 => dff_q_3
        );

    mux_inst_35: MUX2
        port map (
            O => mux_o_35,
            I0 => promx9_inst_16_dout(1),
            I1 => promx9_inst_18_dout(1),
            S0 => dff_q_3
        );

    mux_inst_36: MUX2
        port map (
            O => mux_o_36,
            I0 => mux_o_31,
            I1 => mux_o_32,
            S0 => dff_q_2
        );

    mux_inst_37: MUX2
        port map (
            O => mux_o_37,
            I0 => mux_o_33,
            I1 => mux_o_34,
            S0 => dff_q_2
        );

    mux_inst_39: MUX2
        port map (
            O => mux_o_39,
            I0 => mux_o_36,
            I1 => mux_o_37,
            S0 => dff_q_1
        );

    mux_inst_41: MUX2
        port map (
            O => dout(1),
            I0 => mux_o_39,
            I1 => mux_o_35,
            S0 => dff_q_0
        );

    mux_inst_52: MUX2
        port map (
            O => mux_o_52,
            I0 => promx9_inst_0_dout(2),
            I1 => promx9_inst_1_dout(2),
            S0 => dff_q_3
        );

    mux_inst_53: MUX2
        port map (
            O => mux_o_53,
            I0 => promx9_inst_2_dout(2),
            I1 => promx9_inst_3_dout(2),
            S0 => dff_q_3
        );

    mux_inst_54: MUX2
        port map (
            O => mux_o_54,
            I0 => promx9_inst_4_dout(2),
            I1 => promx9_inst_5_dout(2),
            S0 => dff_q_3
        );

    mux_inst_55: MUX2
        port map (
            O => mux_o_55,
            I0 => promx9_inst_6_dout(2),
            I1 => promx9_inst_7_dout(2),
            S0 => dff_q_3
        );

    mux_inst_56: MUX2
        port map (
            O => mux_o_56,
            I0 => promx9_inst_16_dout(2),
            I1 => promx9_inst_18_dout(2),
            S0 => dff_q_3
        );

    mux_inst_57: MUX2
        port map (
            O => mux_o_57,
            I0 => mux_o_52,
            I1 => mux_o_53,
            S0 => dff_q_2
        );

    mux_inst_58: MUX2
        port map (
            O => mux_o_58,
            I0 => mux_o_54,
            I1 => mux_o_55,
            S0 => dff_q_2
        );

    mux_inst_60: MUX2
        port map (
            O => mux_o_60,
            I0 => mux_o_57,
            I1 => mux_o_58,
            S0 => dff_q_1
        );

    mux_inst_62: MUX2
        port map (
            O => dout(2),
            I0 => mux_o_60,
            I1 => mux_o_56,
            S0 => dff_q_0
        );

    mux_inst_73: MUX2
        port map (
            O => mux_o_73,
            I0 => promx9_inst_0_dout(3),
            I1 => promx9_inst_1_dout(3),
            S0 => dff_q_3
        );

    mux_inst_74: MUX2
        port map (
            O => mux_o_74,
            I0 => promx9_inst_2_dout(3),
            I1 => promx9_inst_3_dout(3),
            S0 => dff_q_3
        );

    mux_inst_75: MUX2
        port map (
            O => mux_o_75,
            I0 => promx9_inst_4_dout(3),
            I1 => promx9_inst_5_dout(3),
            S0 => dff_q_3
        );

    mux_inst_76: MUX2
        port map (
            O => mux_o_76,
            I0 => promx9_inst_6_dout(3),
            I1 => promx9_inst_7_dout(3),
            S0 => dff_q_3
        );

    mux_inst_77: MUX2
        port map (
            O => mux_o_77,
            I0 => promx9_inst_16_dout(3),
            I1 => promx9_inst_18_dout(3),
            S0 => dff_q_3
        );

    mux_inst_78: MUX2
        port map (
            O => mux_o_78,
            I0 => mux_o_73,
            I1 => mux_o_74,
            S0 => dff_q_2
        );

    mux_inst_79: MUX2
        port map (
            O => mux_o_79,
            I0 => mux_o_75,
            I1 => mux_o_76,
            S0 => dff_q_2
        );

    mux_inst_81: MUX2
        port map (
            O => mux_o_81,
            I0 => mux_o_78,
            I1 => mux_o_79,
            S0 => dff_q_1
        );

    mux_inst_83: MUX2
        port map (
            O => dout(3),
            I0 => mux_o_81,
            I1 => mux_o_77,
            S0 => dff_q_0
        );

    mux_inst_94: MUX2
        port map (
            O => mux_o_94,
            I0 => promx9_inst_0_dout(4),
            I1 => promx9_inst_1_dout(4),
            S0 => dff_q_3
        );

    mux_inst_95: MUX2
        port map (
            O => mux_o_95,
            I0 => promx9_inst_2_dout(4),
            I1 => promx9_inst_3_dout(4),
            S0 => dff_q_3
        );

    mux_inst_96: MUX2
        port map (
            O => mux_o_96,
            I0 => promx9_inst_4_dout(4),
            I1 => promx9_inst_5_dout(4),
            S0 => dff_q_3
        );

    mux_inst_97: MUX2
        port map (
            O => mux_o_97,
            I0 => promx9_inst_6_dout(4),
            I1 => promx9_inst_7_dout(4),
            S0 => dff_q_3
        );

    mux_inst_98: MUX2
        port map (
            O => mux_o_98,
            I0 => promx9_inst_16_dout(4),
            I1 => promx9_inst_18_dout(4),
            S0 => dff_q_3
        );

    mux_inst_99: MUX2
        port map (
            O => mux_o_99,
            I0 => mux_o_94,
            I1 => mux_o_95,
            S0 => dff_q_2
        );

    mux_inst_100: MUX2
        port map (
            O => mux_o_100,
            I0 => mux_o_96,
            I1 => mux_o_97,
            S0 => dff_q_2
        );

    mux_inst_102: MUX2
        port map (
            O => mux_o_102,
            I0 => mux_o_99,
            I1 => mux_o_100,
            S0 => dff_q_1
        );

    mux_inst_104: MUX2
        port map (
            O => dout(4),
            I0 => mux_o_102,
            I1 => mux_o_98,
            S0 => dff_q_0
        );

    mux_inst_115: MUX2
        port map (
            O => mux_o_115,
            I0 => promx9_inst_0_dout(5),
            I1 => promx9_inst_1_dout(5),
            S0 => dff_q_3
        );

    mux_inst_116: MUX2
        port map (
            O => mux_o_116,
            I0 => promx9_inst_2_dout(5),
            I1 => promx9_inst_3_dout(5),
            S0 => dff_q_3
        );

    mux_inst_117: MUX2
        port map (
            O => mux_o_117,
            I0 => promx9_inst_4_dout(5),
            I1 => promx9_inst_5_dout(5),
            S0 => dff_q_3
        );

    mux_inst_118: MUX2
        port map (
            O => mux_o_118,
            I0 => promx9_inst_6_dout(5),
            I1 => promx9_inst_7_dout(5),
            S0 => dff_q_3
        );

    mux_inst_119: MUX2
        port map (
            O => mux_o_119,
            I0 => promx9_inst_16_dout(5),
            I1 => promx9_inst_18_dout(5),
            S0 => dff_q_3
        );

    mux_inst_120: MUX2
        port map (
            O => mux_o_120,
            I0 => mux_o_115,
            I1 => mux_o_116,
            S0 => dff_q_2
        );

    mux_inst_121: MUX2
        port map (
            O => mux_o_121,
            I0 => mux_o_117,
            I1 => mux_o_118,
            S0 => dff_q_2
        );

    mux_inst_123: MUX2
        port map (
            O => mux_o_123,
            I0 => mux_o_120,
            I1 => mux_o_121,
            S0 => dff_q_1
        );

    mux_inst_125: MUX2
        port map (
            O => dout(5),
            I0 => mux_o_123,
            I1 => mux_o_119,
            S0 => dff_q_0
        );

    mux_inst_136: MUX2
        port map (
            O => mux_o_136,
            I0 => promx9_inst_0_dout(6),
            I1 => promx9_inst_1_dout(6),
            S0 => dff_q_3
        );

    mux_inst_137: MUX2
        port map (
            O => mux_o_137,
            I0 => promx9_inst_2_dout(6),
            I1 => promx9_inst_3_dout(6),
            S0 => dff_q_3
        );

    mux_inst_138: MUX2
        port map (
            O => mux_o_138,
            I0 => promx9_inst_4_dout(6),
            I1 => promx9_inst_5_dout(6),
            S0 => dff_q_3
        );

    mux_inst_139: MUX2
        port map (
            O => mux_o_139,
            I0 => promx9_inst_6_dout(6),
            I1 => promx9_inst_7_dout(6),
            S0 => dff_q_3
        );

    mux_inst_140: MUX2
        port map (
            O => mux_o_140,
            I0 => promx9_inst_16_dout(6),
            I1 => promx9_inst_18_dout(6),
            S0 => dff_q_3
        );

    mux_inst_141: MUX2
        port map (
            O => mux_o_141,
            I0 => mux_o_136,
            I1 => mux_o_137,
            S0 => dff_q_2
        );

    mux_inst_142: MUX2
        port map (
            O => mux_o_142,
            I0 => mux_o_138,
            I1 => mux_o_139,
            S0 => dff_q_2
        );

    mux_inst_144: MUX2
        port map (
            O => mux_o_144,
            I0 => mux_o_141,
            I1 => mux_o_142,
            S0 => dff_q_1
        );

    mux_inst_146: MUX2
        port map (
            O => dout(6),
            I0 => mux_o_144,
            I1 => mux_o_140,
            S0 => dff_q_0
        );

    mux_inst_157: MUX2
        port map (
            O => mux_o_157,
            I0 => promx9_inst_0_dout(7),
            I1 => promx9_inst_1_dout(7),
            S0 => dff_q_3
        );

    mux_inst_158: MUX2
        port map (
            O => mux_o_158,
            I0 => promx9_inst_2_dout(7),
            I1 => promx9_inst_3_dout(7),
            S0 => dff_q_3
        );

    mux_inst_159: MUX2
        port map (
            O => mux_o_159,
            I0 => promx9_inst_4_dout(7),
            I1 => promx9_inst_5_dout(7),
            S0 => dff_q_3
        );

    mux_inst_160: MUX2
        port map (
            O => mux_o_160,
            I0 => promx9_inst_6_dout(7),
            I1 => promx9_inst_7_dout(7),
            S0 => dff_q_3
        );

    mux_inst_161: MUX2
        port map (
            O => mux_o_161,
            I0 => promx9_inst_16_dout(7),
            I1 => promx9_inst_18_dout(7),
            S0 => dff_q_3
        );

    mux_inst_162: MUX2
        port map (
            O => mux_o_162,
            I0 => mux_o_157,
            I1 => mux_o_158,
            S0 => dff_q_2
        );

    mux_inst_163: MUX2
        port map (
            O => mux_o_163,
            I0 => mux_o_159,
            I1 => mux_o_160,
            S0 => dff_q_2
        );

    mux_inst_165: MUX2
        port map (
            O => mux_o_165,
            I0 => mux_o_162,
            I1 => mux_o_163,
            S0 => dff_q_1
        );

    mux_inst_167: MUX2
        port map (
            O => dout(7),
            I0 => mux_o_165,
            I1 => mux_o_161,
            S0 => dff_q_0
        );

    mux_inst_178: MUX2
        port map (
            O => mux_o_178,
            I0 => promx9_inst_0_dout(8),
            I1 => promx9_inst_1_dout(8),
            S0 => dff_q_3
        );

    mux_inst_179: MUX2
        port map (
            O => mux_o_179,
            I0 => promx9_inst_2_dout(8),
            I1 => promx9_inst_3_dout(8),
            S0 => dff_q_3
        );

    mux_inst_180: MUX2
        port map (
            O => mux_o_180,
            I0 => promx9_inst_4_dout(8),
            I1 => promx9_inst_5_dout(8),
            S0 => dff_q_3
        );

    mux_inst_181: MUX2
        port map (
            O => mux_o_181,
            I0 => promx9_inst_6_dout(8),
            I1 => promx9_inst_7_dout(8),
            S0 => dff_q_3
        );

    mux_inst_182: MUX2
        port map (
            O => mux_o_182,
            I0 => promx9_inst_16_dout(8),
            I1 => promx9_inst_18_dout(8),
            S0 => dff_q_3
        );

    mux_inst_183: MUX2
        port map (
            O => mux_o_183,
            I0 => mux_o_178,
            I1 => mux_o_179,
            S0 => dff_q_2
        );

    mux_inst_184: MUX2
        port map (
            O => mux_o_184,
            I0 => mux_o_180,
            I1 => mux_o_181,
            S0 => dff_q_2
        );

    mux_inst_186: MUX2
        port map (
            O => mux_o_186,
            I0 => mux_o_183,
            I1 => mux_o_184,
            S0 => dff_q_1
        );

    mux_inst_188: MUX2
        port map (
            O => dout(8),
            I0 => mux_o_186,
            I1 => mux_o_182,
            S0 => dff_q_0
        );

    mux_inst_199: MUX2
        port map (
            O => mux_o_199,
            I0 => promx9_inst_8_dout(9),
            I1 => promx9_inst_9_dout(9),
            S0 => dff_q_3
        );

    mux_inst_200: MUX2
        port map (
            O => mux_o_200,
            I0 => promx9_inst_10_dout(9),
            I1 => promx9_inst_11_dout(9),
            S0 => dff_q_3
        );

    mux_inst_201: MUX2
        port map (
            O => mux_o_201,
            I0 => promx9_inst_12_dout(9),
            I1 => promx9_inst_13_dout(9),
            S0 => dff_q_3
        );

    mux_inst_202: MUX2
        port map (
            O => mux_o_202,
            I0 => promx9_inst_14_dout(9),
            I1 => promx9_inst_15_dout(9),
            S0 => dff_q_3
        );

    mux_inst_203: MUX2
        port map (
            O => mux_o_203,
            I0 => promx9_inst_17_dout(9),
            I1 => promx9_inst_18_dout(9),
            S0 => dff_q_3
        );

    mux_inst_204: MUX2
        port map (
            O => mux_o_204,
            I0 => mux_o_199,
            I1 => mux_o_200,
            S0 => dff_q_2
        );

    mux_inst_205: MUX2
        port map (
            O => mux_o_205,
            I0 => mux_o_201,
            I1 => mux_o_202,
            S0 => dff_q_2
        );

    mux_inst_207: MUX2
        port map (
            O => mux_o_207,
            I0 => mux_o_204,
            I1 => mux_o_205,
            S0 => dff_q_1
        );

    mux_inst_209: MUX2
        port map (
            O => dout(9),
            I0 => mux_o_207,
            I1 => mux_o_203,
            S0 => dff_q_0
        );

    mux_inst_220: MUX2
        port map (
            O => mux_o_220,
            I0 => promx9_inst_8_dout(10),
            I1 => promx9_inst_9_dout(10),
            S0 => dff_q_3
        );

    mux_inst_221: MUX2
        port map (
            O => mux_o_221,
            I0 => promx9_inst_10_dout(10),
            I1 => promx9_inst_11_dout(10),
            S0 => dff_q_3
        );

    mux_inst_222: MUX2
        port map (
            O => mux_o_222,
            I0 => promx9_inst_12_dout(10),
            I1 => promx9_inst_13_dout(10),
            S0 => dff_q_3
        );

    mux_inst_223: MUX2
        port map (
            O => mux_o_223,
            I0 => promx9_inst_14_dout(10),
            I1 => promx9_inst_15_dout(10),
            S0 => dff_q_3
        );

    mux_inst_224: MUX2
        port map (
            O => mux_o_224,
            I0 => promx9_inst_17_dout(10),
            I1 => promx9_inst_18_dout(10),
            S0 => dff_q_3
        );

    mux_inst_225: MUX2
        port map (
            O => mux_o_225,
            I0 => mux_o_220,
            I1 => mux_o_221,
            S0 => dff_q_2
        );

    mux_inst_226: MUX2
        port map (
            O => mux_o_226,
            I0 => mux_o_222,
            I1 => mux_o_223,
            S0 => dff_q_2
        );

    mux_inst_228: MUX2
        port map (
            O => mux_o_228,
            I0 => mux_o_225,
            I1 => mux_o_226,
            S0 => dff_q_1
        );

    mux_inst_230: MUX2
        port map (
            O => dout(10),
            I0 => mux_o_228,
            I1 => mux_o_224,
            S0 => dff_q_0
        );

    mux_inst_241: MUX2
        port map (
            O => mux_o_241,
            I0 => promx9_inst_8_dout(11),
            I1 => promx9_inst_9_dout(11),
            S0 => dff_q_3
        );

    mux_inst_242: MUX2
        port map (
            O => mux_o_242,
            I0 => promx9_inst_10_dout(11),
            I1 => promx9_inst_11_dout(11),
            S0 => dff_q_3
        );

    mux_inst_243: MUX2
        port map (
            O => mux_o_243,
            I0 => promx9_inst_12_dout(11),
            I1 => promx9_inst_13_dout(11),
            S0 => dff_q_3
        );

    mux_inst_244: MUX2
        port map (
            O => mux_o_244,
            I0 => promx9_inst_14_dout(11),
            I1 => promx9_inst_15_dout(11),
            S0 => dff_q_3
        );

    mux_inst_245: MUX2
        port map (
            O => mux_o_245,
            I0 => promx9_inst_17_dout(11),
            I1 => promx9_inst_18_dout(11),
            S0 => dff_q_3
        );

    mux_inst_246: MUX2
        port map (
            O => mux_o_246,
            I0 => mux_o_241,
            I1 => mux_o_242,
            S0 => dff_q_2
        );

    mux_inst_247: MUX2
        port map (
            O => mux_o_247,
            I0 => mux_o_243,
            I1 => mux_o_244,
            S0 => dff_q_2
        );

    mux_inst_249: MUX2
        port map (
            O => mux_o_249,
            I0 => mux_o_246,
            I1 => mux_o_247,
            S0 => dff_q_1
        );

    mux_inst_251: MUX2
        port map (
            O => dout(11),
            I0 => mux_o_249,
            I1 => mux_o_245,
            S0 => dff_q_0
        );

    mux_inst_262: MUX2
        port map (
            O => mux_o_262,
            I0 => promx9_inst_8_dout(12),
            I1 => promx9_inst_9_dout(12),
            S0 => dff_q_3
        );

    mux_inst_263: MUX2
        port map (
            O => mux_o_263,
            I0 => promx9_inst_10_dout(12),
            I1 => promx9_inst_11_dout(12),
            S0 => dff_q_3
        );

    mux_inst_264: MUX2
        port map (
            O => mux_o_264,
            I0 => promx9_inst_12_dout(12),
            I1 => promx9_inst_13_dout(12),
            S0 => dff_q_3
        );

    mux_inst_265: MUX2
        port map (
            O => mux_o_265,
            I0 => promx9_inst_14_dout(12),
            I1 => promx9_inst_15_dout(12),
            S0 => dff_q_3
        );

    mux_inst_266: MUX2
        port map (
            O => mux_o_266,
            I0 => promx9_inst_17_dout(12),
            I1 => promx9_inst_18_dout(12),
            S0 => dff_q_3
        );

    mux_inst_267: MUX2
        port map (
            O => mux_o_267,
            I0 => mux_o_262,
            I1 => mux_o_263,
            S0 => dff_q_2
        );

    mux_inst_268: MUX2
        port map (
            O => mux_o_268,
            I0 => mux_o_264,
            I1 => mux_o_265,
            S0 => dff_q_2
        );

    mux_inst_270: MUX2
        port map (
            O => mux_o_270,
            I0 => mux_o_267,
            I1 => mux_o_268,
            S0 => dff_q_1
        );

    mux_inst_272: MUX2
        port map (
            O => dout(12),
            I0 => mux_o_270,
            I1 => mux_o_266,
            S0 => dff_q_0
        );

    mux_inst_283: MUX2
        port map (
            O => mux_o_283,
            I0 => promx9_inst_8_dout(13),
            I1 => promx9_inst_9_dout(13),
            S0 => dff_q_3
        );

    mux_inst_284: MUX2
        port map (
            O => mux_o_284,
            I0 => promx9_inst_10_dout(13),
            I1 => promx9_inst_11_dout(13),
            S0 => dff_q_3
        );

    mux_inst_285: MUX2
        port map (
            O => mux_o_285,
            I0 => promx9_inst_12_dout(13),
            I1 => promx9_inst_13_dout(13),
            S0 => dff_q_3
        );

    mux_inst_286: MUX2
        port map (
            O => mux_o_286,
            I0 => promx9_inst_14_dout(13),
            I1 => promx9_inst_15_dout(13),
            S0 => dff_q_3
        );

    mux_inst_287: MUX2
        port map (
            O => mux_o_287,
            I0 => promx9_inst_17_dout(13),
            I1 => promx9_inst_18_dout(13),
            S0 => dff_q_3
        );

    mux_inst_288: MUX2
        port map (
            O => mux_o_288,
            I0 => mux_o_283,
            I1 => mux_o_284,
            S0 => dff_q_2
        );

    mux_inst_289: MUX2
        port map (
            O => mux_o_289,
            I0 => mux_o_285,
            I1 => mux_o_286,
            S0 => dff_q_2
        );

    mux_inst_291: MUX2
        port map (
            O => mux_o_291,
            I0 => mux_o_288,
            I1 => mux_o_289,
            S0 => dff_q_1
        );

    mux_inst_293: MUX2
        port map (
            O => dout(13),
            I0 => mux_o_291,
            I1 => mux_o_287,
            S0 => dff_q_0
        );

    mux_inst_304: MUX2
        port map (
            O => mux_o_304,
            I0 => promx9_inst_8_dout(14),
            I1 => promx9_inst_9_dout(14),
            S0 => dff_q_3
        );

    mux_inst_305: MUX2
        port map (
            O => mux_o_305,
            I0 => promx9_inst_10_dout(14),
            I1 => promx9_inst_11_dout(14),
            S0 => dff_q_3
        );

    mux_inst_306: MUX2
        port map (
            O => mux_o_306,
            I0 => promx9_inst_12_dout(14),
            I1 => promx9_inst_13_dout(14),
            S0 => dff_q_3
        );

    mux_inst_307: MUX2
        port map (
            O => mux_o_307,
            I0 => promx9_inst_14_dout(14),
            I1 => promx9_inst_15_dout(14),
            S0 => dff_q_3
        );

    mux_inst_308: MUX2
        port map (
            O => mux_o_308,
            I0 => promx9_inst_17_dout(14),
            I1 => promx9_inst_18_dout(14),
            S0 => dff_q_3
        );

    mux_inst_309: MUX2
        port map (
            O => mux_o_309,
            I0 => mux_o_304,
            I1 => mux_o_305,
            S0 => dff_q_2
        );

    mux_inst_310: MUX2
        port map (
            O => mux_o_310,
            I0 => mux_o_306,
            I1 => mux_o_307,
            S0 => dff_q_2
        );

    mux_inst_312: MUX2
        port map (
            O => mux_o_312,
            I0 => mux_o_309,
            I1 => mux_o_310,
            S0 => dff_q_1
        );

    mux_inst_314: MUX2
        port map (
            O => dout(14),
            I0 => mux_o_312,
            I1 => mux_o_308,
            S0 => dff_q_0
        );

    mux_inst_325: MUX2
        port map (
            O => mux_o_325,
            I0 => promx9_inst_8_dout(15),
            I1 => promx9_inst_9_dout(15),
            S0 => dff_q_3
        );

    mux_inst_326: MUX2
        port map (
            O => mux_o_326,
            I0 => promx9_inst_10_dout(15),
            I1 => promx9_inst_11_dout(15),
            S0 => dff_q_3
        );

    mux_inst_327: MUX2
        port map (
            O => mux_o_327,
            I0 => promx9_inst_12_dout(15),
            I1 => promx9_inst_13_dout(15),
            S0 => dff_q_3
        );

    mux_inst_328: MUX2
        port map (
            O => mux_o_328,
            I0 => promx9_inst_14_dout(15),
            I1 => promx9_inst_15_dout(15),
            S0 => dff_q_3
        );

    mux_inst_329: MUX2
        port map (
            O => mux_o_329,
            I0 => promx9_inst_17_dout(15),
            I1 => promx9_inst_18_dout(15),
            S0 => dff_q_3
        );

    mux_inst_330: MUX2
        port map (
            O => mux_o_330,
            I0 => mux_o_325,
            I1 => mux_o_326,
            S0 => dff_q_2
        );

    mux_inst_331: MUX2
        port map (
            O => mux_o_331,
            I0 => mux_o_327,
            I1 => mux_o_328,
            S0 => dff_q_2
        );

    mux_inst_333: MUX2
        port map (
            O => mux_o_333,
            I0 => mux_o_330,
            I1 => mux_o_331,
            S0 => dff_q_1
        );

    mux_inst_335: MUX2
        port map (
            O => dout(15),
            I0 => mux_o_333,
            I1 => mux_o_329,
            S0 => dff_q_0
        );

    mux_inst_346: MUX2
        port map (
            O => mux_o_346,
            I0 => promx9_inst_8_dout(16),
            I1 => promx9_inst_9_dout(16),
            S0 => dff_q_3
        );

    mux_inst_347: MUX2
        port map (
            O => mux_o_347,
            I0 => promx9_inst_10_dout(16),
            I1 => promx9_inst_11_dout(16),
            S0 => dff_q_3
        );

    mux_inst_348: MUX2
        port map (
            O => mux_o_348,
            I0 => promx9_inst_12_dout(16),
            I1 => promx9_inst_13_dout(16),
            S0 => dff_q_3
        );

    mux_inst_349: MUX2
        port map (
            O => mux_o_349,
            I0 => promx9_inst_14_dout(16),
            I1 => promx9_inst_15_dout(16),
            S0 => dff_q_3
        );

    mux_inst_350: MUX2
        port map (
            O => mux_o_350,
            I0 => promx9_inst_17_dout(16),
            I1 => promx9_inst_18_dout(16),
            S0 => dff_q_3
        );

    mux_inst_351: MUX2
        port map (
            O => mux_o_351,
            I0 => mux_o_346,
            I1 => mux_o_347,
            S0 => dff_q_2
        );

    mux_inst_352: MUX2
        port map (
            O => mux_o_352,
            I0 => mux_o_348,
            I1 => mux_o_349,
            S0 => dff_q_2
        );

    mux_inst_354: MUX2
        port map (
            O => mux_o_354,
            I0 => mux_o_351,
            I1 => mux_o_352,
            S0 => dff_q_1
        );

    mux_inst_356: MUX2
        port map (
            O => dout(16),
            I0 => mux_o_354,
            I1 => mux_o_350,
            S0 => dff_q_0
        );

    mux_inst_367: MUX2
        port map (
            O => mux_o_367,
            I0 => promx9_inst_8_dout(17),
            I1 => promx9_inst_9_dout(17),
            S0 => dff_q_3
        );

    mux_inst_368: MUX2
        port map (
            O => mux_o_368,
            I0 => promx9_inst_10_dout(17),
            I1 => promx9_inst_11_dout(17),
            S0 => dff_q_3
        );

    mux_inst_369: MUX2
        port map (
            O => mux_o_369,
            I0 => promx9_inst_12_dout(17),
            I1 => promx9_inst_13_dout(17),
            S0 => dff_q_3
        );

    mux_inst_370: MUX2
        port map (
            O => mux_o_370,
            I0 => promx9_inst_14_dout(17),
            I1 => promx9_inst_15_dout(17),
            S0 => dff_q_3
        );

    mux_inst_371: MUX2
        port map (
            O => mux_o_371,
            I0 => promx9_inst_17_dout(17),
            I1 => promx9_inst_18_dout(17),
            S0 => dff_q_3
        );

    mux_inst_372: MUX2
        port map (
            O => mux_o_372,
            I0 => mux_o_367,
            I1 => mux_o_368,
            S0 => dff_q_2
        );

    mux_inst_373: MUX2
        port map (
            O => mux_o_373,
            I0 => mux_o_369,
            I1 => mux_o_370,
            S0 => dff_q_2
        );

    mux_inst_375: MUX2
        port map (
            O => mux_o_375,
            I0 => mux_o_372,
            I1 => mux_o_373,
            S0 => dff_q_1
        );

    mux_inst_377: MUX2
        port map (
            O => dout(17),
            I0 => mux_o_375,
            I1 => mux_o_371,
            S0 => dff_q_0
        );

end Behavioral; --gato_colorido
