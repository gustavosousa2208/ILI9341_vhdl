--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.07
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Thu Dec 15 15:30:16 2022

library IEEE;
use IEEE.std_logic_1164.all;

entity sprites is
    port (
        dout: out std_logic_vector(1 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(14 downto 0)
    );
end sprites;

architecture Behavioral of sprites is

    signal lut_f_0: std_logic;
    signal lut_f_1: std_logic;
    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_dout: std_logic_vector(0 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout: std_logic_vector(1 downto 1);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout: std_logic_vector(1 downto 0);
    signal dff_q_0: std_logic;
    signal gw_gnd: std_logic;
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);

    -- component declaration
    component LUT2
        generic (
            INIT: in bit_vector := X"0"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic
        );
    end component;

    -- component declaration
    component LUT3
        generic (
            INIT: in bit_vector := X"00"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic
        );
    end component;

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    prom_inst_1_dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    prom_inst_2_dout(1 downto 0) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    lut_inst_0 : LUT2
        generic map (
            INIT => X"2"
        )
        port map (
            F => lut_f_0,
            I0 => ce,
            I1 => ad(14)
        );

    lut_inst_1 : LUT3
        generic map (
            INIT => X"20"
        )
        port map (
            F => lut_f_1,
            I0 => ce,
            I1 => ad(13),
            I2 => ad(14)
        );

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F00FFFF83FC007F9FFF81FF81FF9FFF81F55FFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_01 => X"F83FE3C7FFE007E007F0FFE007E007F87FE0077FF00FC007F0FFF00FE007F8FF",
            INIT_RAM_02 => X"C7E3F807C7E37FE7C3FFC7F03FE3E3C7E3F81FC7E37FE3C7FFC7F07FE1C3C3C3",
            INIT_RAM_03 => X"F07FE3FFF8E7C7E37FFFE3F807F11FE1FFC7FFF8C7C7E3FFFFE3FFC7F13FE3FF",
            INIT_RAM_04 => X"F1C7E0FFF0FFF8FFC7E37EF003E007F1CFF07FE1FFF8FFC7E37EF823F007F18F",
            INIT_RAM_05 => X"C7FFF1E3C7F3FE1FF8FFC7E37EC3C3C7FFF1E3C3FFF83FF8FFC7E37EE003C3C7",
            INIT_RAM_06 => X"C7E3C7E3C003C3E3FF87F8FFC7E37EC7E3C7FFC003C7E3FF0FF8FFC7E37EC7E3",
            INIT_RAM_07 => X"0F7FE007E003F1FFE007E003F8FFE0077EC3C7E3C3F1FFE1C3FFC3F8FFE3C77E",
            INIT_RAM_08 => X"FFFFFFFFF83FF81FF1FFF81FC003F8FFF81FFFF00FF007F1FFF00FC003F8FFF0",
            INIT_RAM_09 => X"1FF81FC003FFFFFFFFFFFBFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0A => X"F7E007E007C007FFFFFFFDFFFFFFF497F00FF00FC0037FFFFFFFFFFFFFFFFFFC",
            INIT_RAM_0B => X"FFFFF7C7E3E3C7F1FF7FAA8BFDF9008FFFFFE3C3E187E3FF7FFFFFFFFFFFFFFF",
            INIT_RAM_0C => X"FFFFFFFFFFC7E3E187F8FFFFFEFFFDFBFFF7FFFFC7E3E3C7F1FFFFFFFFFDFBFF",
            INIT_RAM_0D => X"FFFDFFFFFFE9CFC007F00FFC7FFFFEFFFDFBFFFFFFF7C3C3F00FFC7F7FFFFFFD",
            INIT_RAM_0E => X"7FFEFFFDFFFFFFFFF7C41FC7E3FE3FFFFFFFFDFBFFF7EFFFC00FE3C7FE3F7FFE",
            INIT_RAM_0F => X"FF1F7EFEFFFDFBFBFFFFFFC7FFC7E3FE1F24FEFD83FBFBFFEFF7C7FFC7E3FE3F",
            INIT_RAM_10 => X"E007FF1F7EFEFFFDFBFBFFEFF7E3C7C3C3FF1FFFFEFFFFFBFBFFEFF7C3E7C7E3",
            INIT_RAM_11 => X"FC1FF81FFF9F7EFEFFFFFBFBFFFFFFF00FF00FFF1FFFFEFFFDFBFBFFEA57E007",
            INIT_RAM_12 => X"008FDFDFBFBF007E7EFEFFFFFBFBFFFFFFFFFFFFFFFFFFFFFEFFFDFBFBFFFFFF",
            INIT_RAM_13 => X"FBFFFFFFDFDFFFBFFF7E7EFEFFFFFFFBFFFFFFDFDFFFBFFF7E7EFE8BFD83FBF1",
            INIT_RAM_14 => X"FDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFFFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFF",
            INIT_RAM_15 => X"FEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFFFFFBFFFFFFDFDFFFBFFF7E7EFEFF",
            INIT_RAM_16 => X"FF7FFEFDFDFD009400009FC800007FAA7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7E",
            INIT_RAM_17 => X"FF7FFFFFFEFDFDFFFFF7FFFFDFDFFFFF7FFEFFFEFDFDFFFFF7FFFFDFDFFFFF7F",
            INIT_RAM_18 => X"FFFFFF7FFEFFFEFDFDFFFFFFFFFFDFDFFFFF7FFE7FFEFDFDFFFFFFFFFFFFFFFF",
            INIT_RAM_19 => X"FFFFDFFFFF7FFEFFFEFDFDFFFFFFFFFFDFDFFFFF7FFF7FFEFDFDFFFFF7FFFFFF",
            INIT_RAM_1A => X"FFFFFFDFDFFFFFFFFF7E00FDFD0013F98FFFDFDFD1BF55FE7FFEFDFDFFFFF7FF",
            INIT_RAM_1B => X"FFFFFFFFFFDFDFFFFFFFFE7EFFFDFFFFFBF7FFFFDFDFFFBF7FFF7EFFFDFFFFFB",
            INIT_RAM_1C => X"FDFFFFFFFFFFFFDFDFFFFF7FFE7EFFFDFFFFFBFFFFFFDFDFFFBF7FFF7EFFFDFF",
            INIT_RAM_1D => X"7EFFFDFFFFFBFFFFFFDFDFFFBF7FFE7EFFFDFFFFFBF7FFFFDFDFFFBFFFFF7EFF",
            INIT_RAM_1E => X"FFFE7EFFFDFFFFFFFFFFEFFFDFFFBFFFFF7EFF52000083FFF129BFC8BFBF00AA",
            INIT_RAM_1F => X"BFBFFFFE7EFFFFFFFFFFFFFFFFFFFFFFBFFFFF7EFFFDFFFFFFFFFFEFFFDFBFBF",
            INIT_RAM_20 => X"FFDFBFBFFFFF7EFFFDFFFFFFFFFFEFFFFFFFBFFFFE7EFFFFFFFFFFFFFFFFFFDF",
            INIT_RAM_21 => X"FA9FF01FBFC1007E7EFFFDFFFFFFFFFFEFFFDFBFBFFFFE7EFFFDFFFFFFFFFFFF",
            INIT_RAM_22 => X"FFFFFFEFFFDFFFFFFF7EFFFFFDFFFFFFF7FFFFFFFFFFBFFF7EFE00FDFD0000B7",
            INIT_RAM_23 => X"FDFFFFFFFFFFFFDFFFBFFF7EFEFFFDFFFFFFFFFFFFFFDFFFBFFF7EFFFFFDFDFF",
            INIT_RAM_24 => X"FFFDFDFFFFF7FFEFFFFFFFBFFF7EFEFFFDFFFFFFF7FFFFFFDFFFFFFF7EFFFFFD",
            INIT_RAM_25 => X"107EFEFFFFFFFFFFFFEFFFFFBFFF2110FEFFFDFDFFFFFA5FFFF01FFFFF0070FF",
            INIT_RAM_26 => X"BF21007EFEFFFFFFFFFFFFEFFFFFFFFF21107EFEFFFDFBFFFFFFFFFFFFBFBF21",
            INIT_RAM_27 => X"FFBFFF23087EFEFFFDFFFFFFFFFFFFFFFFBF21087EFEFFFDFBFFFFFFFFFFFFBF",
            INIT_RAM_28 => X"290000BFC100007EFEFFFDFBFFFFFFEFFFFFFFBF230C7EFEFFFFFBFFFFFFEFFF",
            INIT_RAM_29 => X"FFFFFFFFFFFFFF3F037EFFFFFFFBFFFFFFFFFFFFFFFF3F067EFE0083F9000000",
            INIT_RAM_2A => X"FBFFFFFFFFFFFFFFFF0FF07EFFFFFFFFFFFFFFFFFFFFFFFF0FE07EFFFFFFFBFF",
            INIT_RAM_2B => X"FFFFFBFFFFFFFFFFFFFFFF030C7EFFFFFFFFFFFFFFFFFFFFFFFF03087EFFFFFF",
            INIT_RAM_2C => X"7E00000013FBF18FFFC1000000000C7EFFFFFFFBFFFFFFFFFFFFFFFF030C7EFF",
            INIT_RAM_2D => X"FFFEFFFFFDFFFFFBFFFFEFDFFFFFFFFFFF7FFFFDFFFFFBFFFFFFDFFFFFFFFFBE",
            INIT_RAM_2E => X"FFFFFFFF7FFFFDFFFFFBFFFFFFDFFFFFFFFFFE7FFFFFFFFFFFFFFFFFDFFFFFFF",
            INIT_RAM_2F => X"DFFFFFFFFFFF7FFFFDFFFFFBFFFFEFDFFFFFFFFFFEFFFFFFFFFFFFFFFFFFDFFF",
            INIT_RAM_30 => X"FFFFFFFFFFBFFFFE5500FD8BFD13FFF19FDFC1000000AAFFFFFFFFFFFBFFFFFF",
            INIT_RAM_31 => X"FFFFFFFFDFFFFFBFFFFEFFFEFFFDFBFFF7FFFFDFFFFFBFFFFF7FFEFFFDFBFFFF",
            INIT_RAM_32 => X"FDFBFFFFFFFFFFFFFFBFFFFE7FFEFFFDFBFFFFFFFFFFFFFFBFFFFF7FFEFFFDFB",
            INIT_RAM_33 => X"FEFFFDFBFFFFFFFFDFFFFFBFFFFF7FFEFFFDFBFFF7FFFFDFFFFFBFFFFFFFFEFF",
            INIT_RAM_34 => X"7E7FFFFFFFFBFFFFFFFFDFFFFFBF7F7E55FE8BFDFBFD8FFFE92500BFBF00FEFF",
            INIT_RAM_35 => X"BF7F7E7FFFFFFFFBFFFFFFFFDFFFFFFF7F7EFFFFFFFDFBFFF7FFEFDFFFFFBF7F",
            INIT_RAM_36 => X"FFFFBF7F7E7FFFFFFDFBFFFFFFFFDFFFFFFF7F7EFFFFFFFDFBFFFFFFFFDFFFFF",
            INIT_RAM_37 => X"9FDFC100BF7F7EFFFFFFFDFBFFFFFFFFDFFFFFFF7F7EFFFFFFFFFBFFF7FFEFDF",
            INIT_RAM_38 => X"FFFFEFFFDFFFBFFF7E7EFFFDFFFFFFFFFFFFFFDFFFFFFF7E7FFF0083FBFBF900",
            INIT_RAM_39 => X"FFFFFFFFFFFFDFFFBFFF7E7EFFFFFFFBFBFFFFFFFFDFFFFFFF7E7EFFFDFFFBFB",
            INIT_RAM_3A => X"FDFFFBFBFFFFEFFFDFFFFFFF7E7EFFFFFFFFFFFFFFFFFFDFFFBFFF7E7EFFFDFF",
            INIT_RAM_3B => X"7E00FD00A4A4008FF1BFDFBFC1007E7EFFFFFFFBFBFFFFFFFFDFFFBFFF7E7EFF",
            INIT_RAM_3C => X"FFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFF7EFEFFFFFFFFFFFFFFDFFFFFFFFFFE",
            INIT_RAM_3D => X"BFFFFFFF7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFFFFF",
            INIT_RAM_3E => X"DFFFBFFFFFFF7EFEFFFFFFFFFFFFFFDFFFFFFFFFFE7EFEFFFFFFFFFFFFFFDFFF",
            INIT_RAM_3F => X"FFFFFFFFFFFF7FFE7EFE00000083FFF18FDFDFC10000AA7EFEFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F00FFFF83FC007F9FFF81FF81FF9FFF81F55FFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_01 => X"F83FE3C7FFE007E007F0FFE007E007F87FE0077FF00FC007F0FFF00FE007F8FF",
            INIT_RAM_02 => X"C7E3F807C7E37FE7C3FFC7F03FE3E3C7E3F81FC7E37FE3C7FFC7F07FE1C3C3C3",
            INIT_RAM_03 => X"F07FE3FFF8E7C7E37FFFE3F807F11FE1FFC7FFF8C7C7E3FFFFE3FFC7F13FE3FF",
            INIT_RAM_04 => X"F1C7E0FFF0FFF8FFC7E37EF003E007F1CFF07FE1FFF8FFC7E37EF823F007F18F",
            INIT_RAM_05 => X"C7FFF1E3C7F3FE1FF8FFC7E37EC3C3C7FFF1E3C3FFF83FF8FFC7E37EE003C3C7",
            INIT_RAM_06 => X"C7E3C7E3C003C3E3FF87F8FFC7E37EC7E3C7FFC003C7E3FF0FF8FFC7E37EC7E3",
            INIT_RAM_07 => X"0F7FE007E003F1FFE007E003F8FFE0077EC3C7E3C3F1FFE1C3FFC3F8FFE3C77E",
            INIT_RAM_08 => X"FFFFFFFFF83FF81FF1FFF81FC003F8FFF81FFFF00FF007F1FFF00FC003F8FFF0",
            INIT_RAM_09 => X"1FF81FC003FFFFFFFFFFFBFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0A => X"F7E007E007C007FFFFFFFDFFFFFFF497F00FF00FC0037FFFFFFFFFFFFFFFFFFC",
            INIT_RAM_0B => X"FFFFF7C7E3E3C7F1FF7FAA8BFDF9008FFFFFE3C3E187E3FF7FFFFFFFFFFFFFFF",
            INIT_RAM_0C => X"FFFFFFFFFFC7E3E187F8FFFFFEFFFDFBFFF7FFFFC7E3E3C7F1FFFFFFFFFDFBFF",
            INIT_RAM_0D => X"FFFDFFFFFFE9CFC007F00FFC7FFFFEFFFDFBFFFFFFF7C3C3F00FFC7F7FFFFFFD",
            INIT_RAM_0E => X"7FFEFFFDFFFFFFFFF7C41FC7E3FE3FFFFFFFFDFBFFF7EFFFC00FE3C7FE3F7FFE",
            INIT_RAM_0F => X"FF1F7EFEFFFDFBFBFFFFFFC7FFC7E3FE1F24FEFD83FBFBFFEFF7C7FFC7E3FE3F",
            INIT_RAM_10 => X"E007FF1F7EFEFFFDFBFBFFEFF7E3C7C3C3FF1FFFFEFFFFFBFBFFEFF7C3E7C7E3",
            INIT_RAM_11 => X"FC1FF81FFF9F7EFEFFFFFBFBFFFFFFF00FF00FFF1FFFFEFFFDFBFBFFEA57E007",
            INIT_RAM_12 => X"008FDFDFBFBF007E7EFEFFFFFBFBFFFFFFFFFFFFFFFFFFFFFEFFFDFBFBFFFFFF",
            INIT_RAM_13 => X"FBFFFFFFDFDFFFBFFF7E7EFEFFFFFFFBFFFFFFDFDFFFBFFF7E7EFE8BFD83FBF1",
            INIT_RAM_14 => X"FDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFFFFFBFFFFFFDFDFFFBFFF7E7EFEFFFDFF",
            INIT_RAM_15 => X"FEFFFDFFFBFFFFFFDFDFFFBFFF7E7EFEFFFFFFFBFFFFFFDFDFFFBFFF7E7EFEFF",
            INIT_RAM_16 => X"FF7FFEFDFDFD009400009FC800007FAA7EFEFFFDFFFBFFFFFFDFDFFFBFFF7E7E",
            INIT_RAM_17 => X"FF7FFFFFFEFDFDFFFFF7FFFFDFDFFFFF7FFEFFFEFDFDFFFFF7FFFFDFDFFFFF7F",
            INIT_RAM_18 => X"FFFFFF7FFEFFFEFDFDFFFFFFFFFFDFDFFFFF7FFE7FFEFDFDFFFFFFFFFFFFFFFF",
            INIT_RAM_19 => X"FFFFDFFFFF7FFEFFFEFDFDFFFFFFFFFFDFDFFFFF7FFF7FFEFDFDFFFFF7FFFFFF",
            INIT_RAM_1A => X"FFFFFFDFDFFFFFFFFF7E00FDFD0013F98FFFDFDFD1BF55FE7FFEFDFDFFFFF7FF",
            INIT_RAM_1B => X"FFFFFFFFFFDFDFFFFFFFFE7EFFFDFFFFFBF7FFFFDFDFFFBF7FFF7EFFFDFFFFFB",
            INIT_RAM_1C => X"FDFFFFFFFFFFFFDFDFFFFF7FFE7EFFFDFFFFFBFFFFFFDFDFFFBF7FFF7EFFFDFF",
            INIT_RAM_1D => X"7EFFFDFFFFFBFFFFFFDFDFFFBF7FFE7EFFFDFFFFFBF7FFFFDFDFFFBFFFFF7EFF",
            INIT_RAM_1E => X"FFFE7EFFFDFFFFFFFFFFEFFFDFFFBFFFFF7EFF52000083FFF129BFC8BFBF00AA",
            INIT_RAM_1F => X"BFBFFFFE7EFFFFFFFFFFFFFFFFFFFFFFBFFFFF7EFFFDFFFFFFFFFFEFFFDFBFBF",
            INIT_RAM_20 => X"FFDFBFBFFFFF7EFFFDFFFFFFFFFFEFFFFFFFBFFFFE7EFFFFFFFFFFFFFFFFFFDF",
            INIT_RAM_21 => X"FA9FF01FBFC1007E7EFFFDFFFFFFFFFFEFFFDFBFBFFFFE7EFFFDFFFFFFFFFFFF",
            INIT_RAM_22 => X"FFFFFFEFFFDFFFFFFF7EFFFFFDFFFFFFF7FFFFFFFFFFBFFF7EFE00FDFD0000B7",
            INIT_RAM_23 => X"FDFFFFFFFFFFFFDFFFBFFF7EFEFFFDFFFFFFFFFFFFFFDFFFBFFF7EFFFFFDFDFF",
            INIT_RAM_24 => X"FFFDFDFFFFF7FFEFFFFFFFBFFF7EFEFFFDFFFFFFF7FFFFFFDFFFFFFF7EFFFFFD",
            INIT_RAM_25 => X"FF7EFEFFFFFFFFFFFFEFFFFFBFFFFFFFFEFFFDFDFFFFFA5FFFF01FFFFF0C7FFF",
            INIT_RAM_26 => X"BFFFFF7EFEFFFFFFFFFFFFEFFFFFFFFFFFFF7EFEFFFDFBFFFFFFFFFFFFBFBFFF",
            INIT_RAM_27 => X"FFBFFFFFFF7EFEFFFDFFFFFFFFFFFFFFFFBFFFFF7EFEFFFDFBFFFFFFFFFFFFBF",
            INIT_RAM_28 => X"290000BFC1CCFB7EFEFFFDFBFFFFFFEFFFFFFFBFFFFF7EFEFFFFFBFFFFFFEFFF",
            INIT_RAM_29 => X"FFFFFFFFFFFFFFFFFF7EFFFFFFFBFFFFFFFFFFFFFFFFFFFF7EFE0083F9000000",
            INIT_RAM_2A => X"FBFFFFFFFFFFFFFFFFFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFFFFE7EFFFFFFFBFF",
            INIT_RAM_2B => X"FFFFFBFFFFFFFFFFFFFFFFFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFFFFF7EFFFFFF",
            INIT_RAM_2C => X"7E00000013FBF18FFFC10000000CFE7EFFFFFFFBFFFFFFFFFFFFFFFFFFFF7EFF",
            INIT_RAM_2D => X"FFFEFFFFFDFFFFFBFFFFEFDFFFFFFFFFFF7FFFFDFFFFFBFFFFFFDFFFFFFFFFFE",
            INIT_RAM_2E => X"FFFFFFFF7FFFFDFFFFFBFFFFFFDFFFFFFFFFFE7FFFFFFFFFFFFFFFFFDFFFFFFF",
            INIT_RAM_2F => X"DFFFFFFFFFFF7FFFFDFFFFFBFFFFEFDFFFFFFFFFFEFFFFFFFFFFFFFFFFFFDFFF",
            INIT_RAM_30 => X"FFFFFFFFFFBFFFFE5500FD8BFD13FFF19FDFC1000000AAFFFFFFFFFFFBFFFFFF",
            INIT_RAM_31 => X"FFFFFFFFDFFFFFBFFFFEFFFEFFFDFBFFF7FFFFDFFFFFBFFFFF7FFEFFFDFBFFFF",
            INIT_RAM_32 => X"FDFBFFFFFFFFFFFFFFBFFFFE7FFEFFFDFBFFFFFFFFFFFFFFBFFFFF7FFEFFFDFB",
            INIT_RAM_33 => X"FEFFFDFBFFFFFFFFDFFFFFBFFFFF7FFEFFFDFBFFF7FFFFDFFFFFBFFFFFFFFEFF",
            INIT_RAM_34 => X"7E7FFFFFFFFBFFFFFFFFDFFFFFBF7F7E55FE8BFDFBFD8FFFE92500BFBF00FEFF",
            INIT_RAM_35 => X"BF7F7E7FFFFFFFFBFFFFFFFFDFFFFFFF7F7EFFFFFFFDFBFFF7FFEFDFFFFFBF7F",
            INIT_RAM_36 => X"FFFFBF7F7E7FFFFFFDFBFFFFFFFFDFFFFFFF7F7EFFFFFFFDFBFFFFFFFFDFFFFF",
            INIT_RAM_37 => X"9FDFC100BF7F7EFFFFFFFDFBFFFFFFFFDFFFFFFF7F7EFFFFFFFFFBFFF7FFEFDF",
            INIT_RAM_38 => X"FFFFEFFFDFFFBFFF7E7EFFFDFFFFFFFFFFFFFFDFFFFFFF7E7FFF0083FBFBF900",
            INIT_RAM_39 => X"FFFFFFFFFFFFDFFFBFFF7E7EFFFFFFFBFBFFFFFFFFDFFFFFFF7E7EFFFDFFFBFB",
            INIT_RAM_3A => X"FDFFFBFBFFFFEFFFDFFFFFFF7E7EFFFFFFFFFFFFFFFFFFDFFFBFFF7E7EFFFDFF",
            INIT_RAM_3B => X"7E00FD00A4A4008FF1BFDFBFC1007E7EFFFFFFFBFBFFFFFFFFDFFFBFFF7E7EFF",
            INIT_RAM_3C => X"FFFE7EFEFFFFFFFFFFFFFFDFFFBFFFFFFF7EFEFFFFFFFFFFFFFFDFFFFFFFFFFE",
            INIT_RAM_3D => X"BFFFFFFF7EFEFFFFFFFFFFFFFFDFFFBFFFFFFE7EFEFFFFFFFFFFFFFFDFFFFFFF",
            INIT_RAM_3E => X"DFFFBFFFFFFF7EFEFFFFFFFFFFFFFFDFFFFFFFFFFE7EFEFFFFFFFFFFFFFFDFFF",
            INIT_RAM_3F => X"FFFFFFFFFFFF7FFE7EFE00000083FFF18FDFDFC10000AA7EFEFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_0,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"FFFFFFFFFCFFFFFFF3FFCFFFFFFF3FFFFFFF3FFFFFFCFFFFFFF3FFFFFFCFFFFF",
            INIT_RAM_01 => X"FFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFCFFFFFFFFFFFFFFF3FFFFFFCF",
            INIT_RAM_02 => X"FFFFFFCFFFFFFFFFFFFFFFFFF3FFCFFFFFFF3FFFFFFF3FFFFFFCFFFFFFF3FFFF",
            INIT_RAM_03 => X"FFF3FFFFFFCFFFFFFFFFFFFFFFFFFFFFCFFFFFFF3FFFFFFCFFFFFFFCFFFFFFF3",
            INIT_RAM_04 => X"FFFFFFF3FFFFFFCFFFFFFFFFFCFFFFFFF3FFFFFFFFFF3FFFFFFF3FFFFFFFFFFF",
            INIT_RAM_05 => X"FFFFFFFFFFF3FFFFFFCFFFFFFFFFFFFFFFFFF3FFCFFFFFFF3FFFFFFFFFFFFFFC",
            INIT_RAM_06 => X"3FFFCCCCFFF3FFF3FFCFFFCFFFFFFFFFFF030000C3FFF003CFFF3FFFFFFCFFFF",
            INIT_RAM_07 => X"3FFC3FFCFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFCFFFFFFF3FFF3FFC",
            INIT_RAM_08 => X"3FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFFFFFFFFFCFFFFFFFFFFCFFFFFFF3FFF",
            INIT_RAM_09 => X"FFFF3FFF3FFC3FFCFFFFFFFFFFFFFFCFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0A => X"FFFFFFFF3FFF3FFC3FFCFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF",
            INIT_RAM_0B => X"FFFFCFFFFFFF3FFF3FFC3FFCFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_0C => X"FFFFFFFFFFFFFFFF3FFF3FFC3FFCFFFFFFFFFFFFFFCFFFFFFF3FFFFFFCFFFFFF",
            INIT_RAM_0D => X"C3FFF3FFF003CFFFF3033FFF3FFC3FFCFFFFFFF3FFFFFFCFFFFFFF3FFFFFFFFF",
            INIT_RAM_0E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFC3FFCFFFFC00FFFF3CC300000C3300000",
            INIT_RAM_0F => X"FFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFF3FFCFFFFFFF3FFFFFFFFFFFFFFFF",
            INIT_RAM_10 => X"FFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFCFFFFFFFFFFF3FFFFFFFFFFFF",
            INIT_RAM_11 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFCFFFFFFF3FFFFFFFF",
            INIT_RAM_12 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFCFFFFFFFFFFFFFFFF",
            INIT_RAM_13 => X"FFF3FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFF3FFCFFFFFFFF",
            INIT_RAM_14 => X"FFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFF3FFCFFFFFFFF",
            INIT_RAM_15 => X"0C300000330C0000000000000000000000000C3300000000000000000C303FFC"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ad(14),
            CLK => clk,
            CE => ce
        );

    mux_inst_2: MUX2
        port map (
            O => dout(0),
            I0 => prom_inst_0_dout(0),
            I1 => prom_inst_2_dout(0),
            S0 => dff_q_0
        );

    mux_inst_5: MUX2
        port map (
            O => dout(1),
            I0 => prom_inst_1_dout(1),
            I1 => prom_inst_2_dout(1),
            S0 => dff_q_0
        );

end Behavioral; --sprites
