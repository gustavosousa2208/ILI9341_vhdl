//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Mon Dec 12 22:06:27 2022

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [1:0] douta;
output [1:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [14:0] ada;
input [1:0] dina;
input [14:0] adb;
input [1:0] dinb;

wire [14:0] dpb_inst_0_douta_w;
wire [0:0] dpb_inst_0_douta;
wire [14:0] dpb_inst_0_doutb_w;
wire [0:0] dpb_inst_0_doutb;
wire [14:0] dpb_inst_1_douta_w;
wire [1:1] dpb_inst_1_douta;
wire [14:0] dpb_inst_1_doutb_w;
wire [1:1] dpb_inst_1_doutb;
wire [13:0] dpb_inst_2_douta_w;
wire [1:0] dpb_inst_2_douta;
wire [13:0] dpb_inst_2_doutb_w;
wire [1:0] dpb_inst_2_doutb;
wire dff_q_0;
wire dff_q_1;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[14:0],dpb_inst_0_douta[0]}),
    .DOB({dpb_inst_0_doutb_w[14:0],dpb_inst_0_doutb[0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[0]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 1;
defparam dpb_inst_0.BIT_WIDTH_1 = 1;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFEFFFFFFFE00000000000000000000FE000000000000000000;
defparam dpb_inst_0.INIT_RAM_01 = 256'hFFFFFFFE7FFFFFFFFFFF7F7FFFFFFFFFFFFFFFFEFFFFFFFE7FFFFFFFFFFF7F7F;
defparam dpb_inst_0.INIT_RAM_02 = 256'hFFFF7F7FFFFFFFFFFFFFFFFEFFFFFFFE7FFFFFFFFFFF7F7FFFFFFFFFFFFFFFFE;
defparam dpb_inst_0.INIT_RAM_03 = 256'hFFFFFFFEFFFFFFFE7FFFFFFFFFFF7F7FFFFFFFFFFFFFFFFEFFFFFFFE7FFFFFFF;
defparam dpb_inst_0.INIT_RAM_04 = 256'h00007F00007F7F7F0000000000FE0000FEFE00FE7FFFFFFFFFFF7F7FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_05 = 256'h7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE;
defparam dpb_inst_0.INIT_RAM_06 = 256'hFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F;
defparam dpb_inst_0.INIT_RAM_07 = 256'h7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFF;
defparam dpb_inst_0.INIT_RAM_08 = 256'hFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF;
defparam dpb_inst_0.INIT_RAM_09 = 256'h7F7F00007F7F007F7F00FEFEFE00000000FEFE007FFF7FFF7FFFFF7F7FFFFEFF;
defparam dpb_inst_0.INIT_RAM_0A = 256'h7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE;
defparam dpb_inst_0.INIT_RAM_0B = 256'hFEFEFFFE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7FFF7F7FFF;
defparam dpb_inst_0.INIT_RAM_0C = 256'hFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFF;
defparam dpb_inst_0.INIT_RAM_0D = 256'h0000FEFEFEFE00FE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7F;
defparam dpb_inst_0.INIT_RAM_0E = 256'h7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE00007F7F007F7F007F7F0000;
defparam dpb_inst_0.INIT_RAM_0F = 256'h7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE;
defparam dpb_inst_0.INIT_RAM_10 = 256'hFFFEFFFE7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F7F7FFF7F;
defparam dpb_inst_0.INIT_RAM_11 = 256'h7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFE;
defparam dpb_inst_0.INIT_RAM_12 = 256'hFE0000000000FE007FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F;
defparam dpb_inst_0.INIT_RAM_13 = 256'h7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE7F7F007F7F00007F7F0000FE;
defparam dpb_inst_0.INIT_RAM_14 = 256'h7FFFFEFEFEFFFEFFFFFFFEFE7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE;
defparam dpb_inst_0.INIT_RAM_15 = 256'hFFFFFEFE7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE7F7FFF7F7FFFFFFF;
defparam dpb_inst_0.INIT_RAM_16 = 256'h7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFF;
defparam dpb_inst_0.INIT_RAM_17 = 256'hFEFEFFFFFEFFFFFE7F007F7F0000007F0000FEFEFEFEFE0000FE00FE7F7FFF7F;
defparam dpb_inst_0.INIT_RAM_18 = 256'h7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFE;
defparam dpb_inst_0.INIT_RAM_19 = 256'hFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE;
defparam dpb_inst_0.INIT_RAM_1A = 256'hFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7F;
defparam dpb_inst_0.INIT_RAM_1B = 256'h7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFF;
defparam dpb_inst_0.INIT_RAM_1C = 256'hFFFEFFFFFEFFFEFE7F7F007F007F7F007F7FFEFE00FE0000FE00FE007F7FFF7F;
defparam dpb_inst_0.INIT_RAM_1D = 256'h7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFFFEFFFEFE7F7FFFFF7FFF7FFFFF7FFEFF;
defparam dpb_inst_0.INIT_RAM_1E = 256'hFF7FFEFFFFFEFFFFFEFFFEFE7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFFFEFFFEFE;
defparam dpb_inst_0.INIT_RAM_1F = 256'hFEFFFEFE7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFFFEFFFEFE7F7FFFFF7FFF7FFF;
defparam dpb_inst_0.INIT_RAM_20 = 256'h7F0000007F7F00000000FE0000FE00FE7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFF;
defparam dpb_inst_0.INIT_RAM_21 = 256'hFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE7F00007F;
defparam dpb_inst_0.INIT_RAM_22 = 256'h7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFF;
defparam dpb_inst_0.INIT_RAM_23 = 256'h7F7F7FFFFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE;
defparam dpb_inst_0.INIT_RAM_24 = 256'hFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF;
defparam dpb_inst_0.INIT_RAM_25 = 256'hFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFF;
defparam dpb_inst_0.INIT_RAM_26 = 256'hFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7F007F;
defparam dpb_inst_0.INIT_RAM_27 = 256'h7F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7FFF7FFEFE;
defparam dpb_inst_0.INIT_RAM_28 = 256'hFF7FFEFEFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE;
defparam dpb_inst_0.INIT_RAM_29 = 256'h00FE00007F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7F;
defparam dpb_inst_0.INIT_RAM_2A = 256'h7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE7F00007F00007F000000000000FEFE00;
defparam dpb_inst_0.INIT_RAM_2B = 256'hFFFEFFFEFFFEFFFE7FFF7FFF7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE7FFF7FFF;
defparam dpb_inst_0.INIT_RAM_2C = 256'h7FFF7FFF7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE7FFF7FFF7FFF7FFFFF7FFFFE;
defparam dpb_inst_0.INIT_RAM_2D = 256'hFF7FFFFEFFFEFFFEFFFEFFFE7FFF7FFF7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE;
defparam dpb_inst_0.INIT_RAM_2E = 256'hFFFEFFFE007F7F007F0000007F7F7EFE000000FEFE0000FE7FFF7FFF7FFF7FFF;
defparam dpb_inst_0.INIT_RAM_2F = 256'hFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFE;
defparam dpb_inst_0.INIT_RAM_30 = 256'hFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFF;
defparam dpb_inst_0.INIT_RAM_31 = 256'h7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFF;
defparam dpb_inst_0.INIT_RAM_32 = 256'h7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE;
defparam dpb_inst_0.INIT_RAM_33 = 256'hFEFEFEFE7F7F007F007F7F7F7F7F000000000000FEFEFE007FFF7FFFFFFF7FFF;
defparam dpb_inst_0.INIT_RAM_34 = 256'hFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFF;
defparam dpb_inst_0.INIT_RAM_35 = 256'hFFFEFFFFFEFEFEFE7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE7F7FFFFF;
defparam dpb_inst_0.INIT_RAM_36 = 256'h7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE7F7FFFFFFF7F7F7F7F7FFFFE;
defparam dpb_inst_0.INIT_RAM_37 = 256'h7F00FE00FEFEFE0000FEFEFE7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE;
defparam dpb_inst_0.INIT_RAM_38 = 256'hFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7F0000007F7F7F7F;
defparam dpb_inst_0.INIT_RAM_39 = 256'hFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFE;
defparam dpb_inst_0.INIT_RAM_3A = 256'hFEFEFFFEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7FFF7F7F;
defparam dpb_inst_0.INIT_RAM_3B = 256'h7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFF;
defparam dpb_inst_0.INIT_RAM_3C = 256'h7F00000000FE00FEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE;
defparam dpb_inst_0.INIT_RAM_3D = 256'hFEFFFEFE7F7FFF7F7FFFFF7F7F7FFEFFFFFEFFFEFEFFFEFE7F7F7F7F0000007F;
defparam dpb_inst_0.INIT_RAM_3E = 256'h7FFFFF7F7F7FFEFFFFFEFFFEFEFFFEFE7F7FFF7F7FFFFF7F7F7FFEFFFFFEFFFE;
defparam dpb_inst_0.INIT_RAM_3F = 256'hFFFEFFFEFEFFFEFE7F7FFF7F7FFFFF7F7F7FFEFFFFFEFFFEFEFFFEFE7F7FFF7F;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[14:0],dpb_inst_1_douta[1]}),
    .DOB({dpb_inst_1_doutb_w[14:0],dpb_inst_1_doutb[1]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 1;
defparam dpb_inst_1.BIT_WIDTH_1 = 1;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFEFFFFFFFE00000000000000000000FE000000000000000000;
defparam dpb_inst_1.INIT_RAM_01 = 256'hFFFFFFFE7FFFFFFFFFFF7F7FFFFFFFFFFFFFFFFEFFFFFFFE7FFFFFFFFFFF7F7F;
defparam dpb_inst_1.INIT_RAM_02 = 256'hFFFF7F7FFFFFFFFFFFFFFFFEFFFFFFFE7FFFFFFFFFFF7F7FFFFFFFFFFFFFFFFE;
defparam dpb_inst_1.INIT_RAM_03 = 256'hFFFFFFFEFFFFFFFE7FFFFFFFFFFF7F7FFFFFFFFFFFFFFFFEFFFFFFFE7FFFFFFF;
defparam dpb_inst_1.INIT_RAM_04 = 256'h00007F00007F7F7F0000000000FE0000FEFE00FE7FFFFFFFFFFF7F7FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_05 = 256'h7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE;
defparam dpb_inst_1.INIT_RAM_06 = 256'hFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F;
defparam dpb_inst_1.INIT_RAM_07 = 256'h7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFF;
defparam dpb_inst_1.INIT_RAM_08 = 256'hFEFFFFFFFEFFFEFE7FFF7FFF7FFFFF7F7FFFFEFFFEFFFFFFFEFFFEFE7FFF7FFF;
defparam dpb_inst_1.INIT_RAM_09 = 256'h7F7F00007F7F007F7F00FEFEFE00000000FEFE007FFF7FFF7FFFFF7F7FFFFEFF;
defparam dpb_inst_1.INIT_RAM_0A = 256'h7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE;
defparam dpb_inst_1.INIT_RAM_0B = 256'hFEFEFFFE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7FFF7F7FFF;
defparam dpb_inst_1.INIT_RAM_0C = 256'hFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFF;
defparam dpb_inst_1.INIT_RAM_0D = 256'h0000FEFEFEFE00FE7F7FFF7FFF7F7FFF7F7FFFFEFFFFFEFFFEFEFFFE7F7FFF7F;
defparam dpb_inst_1.INIT_RAM_0E = 256'h7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE00007F7F007F7F007F7F0000;
defparam dpb_inst_1.INIT_RAM_0F = 256'h7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE;
defparam dpb_inst_1.INIT_RAM_10 = 256'hFFFEFFFE7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F7F7FFF7F;
defparam dpb_inst_1.INIT_RAM_11 = 256'h7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFE;
defparam dpb_inst_1.INIT_RAM_12 = 256'hFE0000000000FE007FFFFF7F7F7FFF7F7F7FFFFEFFFFFFFEFFFEFFFE7FFFFF7F;
defparam dpb_inst_1.INIT_RAM_13 = 256'h7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE7F7F007F7F00007F7F0000FE;
defparam dpb_inst_1.INIT_RAM_14 = 256'h7FFFFEFEFEFFFEFFFFFFFEFE7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE;
defparam dpb_inst_1.INIT_RAM_15 = 256'hFFFFFEFE7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE7F7FFF7F7FFFFFFF;
defparam dpb_inst_1.INIT_RAM_16 = 256'h7FFFFFFF7FFFFEFEFEFFFEFFFFFFFEFE7F7FFF7F7FFFFFFF7FFFFEFEFEFFFEFF;
defparam dpb_inst_1.INIT_RAM_17 = 256'hFEFEFFFFFEFFFFFE7F007F7F0000007F0000FEFEFEFEFE0000FE00FE7F7FFF7F;
defparam dpb_inst_1.INIT_RAM_18 = 256'h7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFE;
defparam dpb_inst_1.INIT_RAM_19 = 256'hFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE;
defparam dpb_inst_1.INIT_RAM_1A = 256'hFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7F;
defparam dpb_inst_1.INIT_RAM_1B = 256'h7FFFFF7FFF7FFEFEFEFEFFFFFEFFFFFE7F7FFF7F7FFFFF7FFF7FFEFEFEFEFFFF;
defparam dpb_inst_1.INIT_RAM_1C = 256'hFFFEFFFFFEFFFEFE7F7F007F007F7F007F7FFEFE00FE0000FE00FE007F7FFF7F;
defparam dpb_inst_1.INIT_RAM_1D = 256'h7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFFFEFFFEFE7F7FFFFF7FFF7FFFFF7FFEFF;
defparam dpb_inst_1.INIT_RAM_1E = 256'hFF7FFEFFFFFEFFFFFEFFFEFE7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFFFEFFFEFE;
defparam dpb_inst_1.INIT_RAM_1F = 256'hFEFFFEFE7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFFFEFFFEFE7F7FFFFF7FFF7FFF;
defparam dpb_inst_1.INIT_RAM_20 = 256'h7F0000007F7F00000000FE0000FE00FE7F7FFFFF7FFF7FFFFF7FFEFFFFFEFFFF;
defparam dpb_inst_1.INIT_RAM_21 = 256'hFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE7F00007F;
defparam dpb_inst_1.INIT_RAM_22 = 256'h7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFF;
defparam dpb_inst_1.INIT_RAM_23 = 256'h7F7F7FFFFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE;
defparam dpb_inst_1.INIT_RAM_24 = 256'hFFFEFEFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFFFFFEFEFE7F7FFFFF7F7FFFFF;
defparam dpb_inst_1.INIT_RAM_25 = 256'hFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7FFFFF7F7FFFFF7F7F7FFFFEFEFEFF;
defparam dpb_inst_1.INIT_RAM_26 = 256'hFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7F007F;
defparam dpb_inst_1.INIT_RAM_27 = 256'h7F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7FFF7FFEFE;
defparam dpb_inst_1.INIT_RAM_28 = 256'hFF7FFEFEFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE;
defparam dpb_inst_1.INIT_RAM_29 = 256'h00FE00007F7FFF7FFF7FFF7FFF7FFEFEFFFEFEFFFEFFFFFE7F7FFF7FFF7FFF7F;
defparam dpb_inst_1.INIT_RAM_2A = 256'h7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE7F00007F00007F000000000000FEFE00;
defparam dpb_inst_1.INIT_RAM_2B = 256'hFFFEFFFEFFFEFFFE7FFF7FFF7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE7FFF7FFF;
defparam dpb_inst_1.INIT_RAM_2C = 256'h7FFF7FFF7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE7FFF7FFF7FFF7FFFFF7FFFFE;
defparam dpb_inst_1.INIT_RAM_2D = 256'hFF7FFFFEFFFEFFFEFFFEFFFE7FFF7FFF7FFF7FFFFF7FFFFEFFFEFFFEFFFEFFFE;
defparam dpb_inst_1.INIT_RAM_2E = 256'hFFFEFFFE007F7F007F0000007F7F7EFE000000FEFE0000FE7FFF7FFF7FFF7FFF;
defparam dpb_inst_1.INIT_RAM_2F = 256'hFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFE;
defparam dpb_inst_1.INIT_RAM_30 = 256'hFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFF;
defparam dpb_inst_1.INIT_RAM_31 = 256'h7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFF;
defparam dpb_inst_1.INIT_RAM_32 = 256'h7F7F7EFFFFFFFFFEFFFEFFFE7FFF7FFFFFFF7FFF7F7F7EFFFFFFFFFEFFFEFFFE;
defparam dpb_inst_1.INIT_RAM_33 = 256'hFEFEFEFE7F7F007F007F7F7F7F7F000000000000FEFEFE007FFF7FFFFFFF7FFF;
defparam dpb_inst_1.INIT_RAM_34 = 256'hFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFF;
defparam dpb_inst_1.INIT_RAM_35 = 256'hFFFEFFFFFEFEFEFE7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE7F7FFFFF;
defparam dpb_inst_1.INIT_RAM_36 = 256'h7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE7F7FFFFFFF7F7F7F7F7FFFFE;
defparam dpb_inst_1.INIT_RAM_37 = 256'h7F00FE00FEFEFE0000FEFEFE7F7FFFFFFF7F7F7F7F7FFFFEFFFEFFFFFEFEFEFE;
defparam dpb_inst_1.INIT_RAM_38 = 256'hFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7F0000007F7F7F7F;
defparam dpb_inst_1.INIT_RAM_39 = 256'hFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFE;
defparam dpb_inst_1.INIT_RAM_3A = 256'hFEFEFFFEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7FFF7F7F;
defparam dpb_inst_1.INIT_RAM_3B = 256'h7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFF;
defparam dpb_inst_1.INIT_RAM_3C = 256'h7F00000000FE00FEFEFEFEFE7FFF7F7FFF7FFF7F7FFFFFFFFEFEFFFEFEFEFEFE;
defparam dpb_inst_1.INIT_RAM_3D = 256'hFEFFFEFE7F7FFF7F7FFFFF7F7F7FFEFFFFFEFFFEFEFFFEFE7F7F7F7F0000007F;
defparam dpb_inst_1.INIT_RAM_3E = 256'h7FFFFF7F7F7FFEFFFFFEFFFEFEFFFEFE7F7FFF7F7FFFFF7F7F7FFEFFFFFEFFFE;
defparam dpb_inst_1.INIT_RAM_3F = 256'hFFFEFFFEFEFFFEFE7F7FFF7F7FFFFF7F7F7FFEFFFFFEFFFEFEFFFEFE7F7FFF7F;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[13:0],dpb_inst_2_douta[1:0]}),
    .DOB({dpb_inst_2_doutb_w[13:0],dpb_inst_2_doutb[1:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1:0]}),
    .ADB({adb[12:0],gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1:0]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b0;
defparam dpb_inst_2.READ_MODE1 = 1'b0;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 2;
defparam dpb_inst_2.BIT_WIDTH_1 = 2;
defparam dpb_inst_2.BLK_SEL_0 = 3'b010;
defparam dpb_inst_2.BLK_SEL_1 = 3'b010;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'hFFFCFFFFFFFCFFFC3FFF3FFFFFFF3FFF3FFFFFFFFFFF3FFF3FFF3FFFFFFCFFFF;
defparam dpb_inst_2.INIT_RAM_01 = 256'h3FFF3FFFFFFF3FFF3FFFFFFFFFFF3FFF3FFF3FFFFFFCFFFFFFFFFFFCFFFFFFFC;
defparam dpb_inst_2.INIT_RAM_02 = 256'h3FFF00003FFF3FFF3FFF3FFF3FFCFFFC00000000FFFC0000FFFCFFFC0000FFFC;
defparam dpb_inst_2.INIT_RAM_03 = 256'h3FFF3FFF3FFCFFFCFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFC3FFF000000003FFF;
defparam dpb_inst_2.INIT_RAM_04 = 256'hFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFC3FFFFFFFFFFF3FFF3FFFFFFF3FFF3FFF;
defparam dpb_inst_2.INIT_RAM_05 = 256'hFFFCFFFFFFFFFFFC3FFFFFFFFFFF3FFF3FFFFFFF3FFF3FFF3FFF3FFF3FFCFFFC;
defparam dpb_inst_2.INIT_RAM_06 = 256'h3FFFFFFFFFFF3FFF3FFFFFFF3FFF3FFF3FFF3FFF3FFCFFFCFFFCFFFFFFFCFFFF;
defparam dpb_inst_2.INIT_RAM_07 = 256'h3FFFFFFF3FFF3FFF3FFF3FFF3FFCFFFCFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFC;
defparam dpb_inst_2.INIT_RAM_08 = 256'h3FFF3FFF3FFCFFFCFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFC3FFFFFFFFFFF3FFF;
defparam dpb_inst_2.INIT_RAM_09 = 256'hFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFC3FFFFFFFFFFF3FFF3FFFFFFF3FFF3FFF;
defparam dpb_inst_2.INIT_RAM_0A = 256'hFFFCFFFFFFFFFFFC3FFFFFFFFFFF3FFF3FFFFFFF3FFF3FFF3FFF3FFF3FFCFFFC;
defparam dpb_inst_2.INIT_RAM_0B = 256'h3FFFFFFFFFFF3FFF3FFFFFFF3FFF3FFF3FFF3FFF3FFCFFFCFFFCFFFFFFFCFFFF;
defparam dpb_inst_2.INIT_RAM_0C = 256'h000000003FFF3FFF3FFF3FFF0000FFFCFFFCFFFC0000FFFCFFFC00000000FFFC;
defparam dpb_inst_2.INIT_RAM_0D = 256'hFFFF3FFFFFFFFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFFFFFC000000003FFF3FFF;
defparam dpb_inst_2.INIT_RAM_0E = 256'hFFFFFFFCFFFFFFFCFFFFFFFFFFFFFFFC3FFFFFFFFFFF3FFFFFFFFFFFFFFF3FFF;
defparam dpb_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFC3FFFFFFFFFFF3FFFFFFFFFFFFFFF3FFFFFFF3FFFFFFFFFFC;
defparam dpb_inst_2.INIT_RAM_10 = 256'h3FFFFFFFFFFF3FFFFFFFFFFFFFFF3FFFFFFF3FFFFFFFFFFCFFFFFFFCFFFFFFFC;
defparam dpb_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFF3FFFFFFF3FFFFFFFFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFFFFFC;
defparam dpb_inst_2.INIT_RAM_12 = 256'hFFFF3FFFFFFFFFFCFFFFFFFCFFFFFFFCFFFFFFFFFFFFFFFC3FFFFFFFFFFF3FFF;
defparam dpb_inst_2.INIT_RAM_13 = 256'hFFFFFFFCFFFFFFFCFFFFFFFFFFFFFFFC3FFFFFFFFFFF3FFFFFFFFFFFFFFF3FFF;
defparam dpb_inst_2.INIT_RAM_14 = 256'h00000000000000003FFFFFFFFFFF3FFFFFFFFFFFFFFF3FFFFFFF3FFFFFFFFFFC;
defparam dpb_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000003FFF000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[14]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb_w)
);
MUX2 mux_inst_2 (
  .O(douta[0]),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_2_douta[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(douta[1]),
  .I0(dpb_inst_1_douta[1]),
  .I1(dpb_inst_2_douta[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(doutb[0]),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_2_doutb[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_11 (
  .O(doutb[1]),
  .I0(dpb_inst_1_doutb[1]),
  .I1(dpb_inst_2_doutb[1]),
  .S0(dff_q_1)
);
endmodule //Gowin_DPB
