--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.07
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Thu Dec 15 12:09:20 2022

library IEEE;
use IEEE.std_logic_1164.all;

entity gato_colorido is
    port (
        dout: out std_logic_vector(17 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(14 downto 0)
    );
end gato_colorido;

architecture Behavioral of gato_colorido is

    signal lut_f_0: std_logic;
    signal lut_f_1: std_logic;
    signal lut_f_2: std_logic;
    signal lut_f_3: std_logic;
    signal lut_f_4: std_logic;
    signal lut_f_5: std_logic;
    signal lut_f_6: std_logic;
    signal lut_f_7: std_logic;
    signal lut_f_8: std_logic;
    signal lut_f_9: std_logic;
    signal lut_f_10: std_logic;
    signal lut_f_11: std_logic;
    signal lut_f_12: std_logic;
    signal lut_f_13: std_logic;
    signal lut_f_14: std_logic;
    signal lut_f_15: std_logic;
    signal lut_f_16: std_logic;
    signal lut_f_17: std_logic;
    signal lut_f_18: std_logic;
    signal lut_f_19: std_logic;
    signal promx9_inst_0_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_0_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_1_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_1_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_2_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_2_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_3_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_3_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_4_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_4_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_5_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_5_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_6_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_6_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_7_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_7_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_8_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_8_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_9_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_9_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_10_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_10_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_11_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_11_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_12_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_12_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_13_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_13_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_14_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_14_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_15_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_15_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_16_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_16_dout: std_logic_vector(8 downto 0);
    signal promx9_inst_17_dout_w: std_logic_vector(26 downto 0);
    signal promx9_inst_17_dout: std_logic_vector(17 downto 9);
    signal promx9_inst_18_dout_w: std_logic_vector(17 downto 0);
    signal promx9_inst_18_dout: std_logic_vector(17 downto 0);
    signal dff_q_0: std_logic;
    signal dff_q_1: std_logic;
    signal dff_q_2: std_logic;
    signal dff_q_3: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_11: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_13: std_logic;
    signal mux_o_14: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_31: std_logic;
    signal mux_o_32: std_logic;
    signal mux_o_33: std_logic;
    signal mux_o_34: std_logic;
    signal mux_o_35: std_logic;
    signal mux_o_36: std_logic;
    signal mux_o_37: std_logic;
    signal mux_o_39: std_logic;
    signal mux_o_52: std_logic;
    signal mux_o_53: std_logic;
    signal mux_o_54: std_logic;
    signal mux_o_55: std_logic;
    signal mux_o_56: std_logic;
    signal mux_o_57: std_logic;
    signal mux_o_58: std_logic;
    signal mux_o_60: std_logic;
    signal mux_o_73: std_logic;
    signal mux_o_74: std_logic;
    signal mux_o_75: std_logic;
    signal mux_o_76: std_logic;
    signal mux_o_77: std_logic;
    signal mux_o_78: std_logic;
    signal mux_o_79: std_logic;
    signal mux_o_81: std_logic;
    signal mux_o_94: std_logic;
    signal mux_o_95: std_logic;
    signal mux_o_96: std_logic;
    signal mux_o_97: std_logic;
    signal mux_o_98: std_logic;
    signal mux_o_99: std_logic;
    signal mux_o_100: std_logic;
    signal mux_o_102: std_logic;
    signal mux_o_115: std_logic;
    signal mux_o_116: std_logic;
    signal mux_o_117: std_logic;
    signal mux_o_118: std_logic;
    signal mux_o_119: std_logic;
    signal mux_o_120: std_logic;
    signal mux_o_121: std_logic;
    signal mux_o_123: std_logic;
    signal mux_o_136: std_logic;
    signal mux_o_137: std_logic;
    signal mux_o_138: std_logic;
    signal mux_o_139: std_logic;
    signal mux_o_140: std_logic;
    signal mux_o_141: std_logic;
    signal mux_o_142: std_logic;
    signal mux_o_144: std_logic;
    signal mux_o_157: std_logic;
    signal mux_o_158: std_logic;
    signal mux_o_159: std_logic;
    signal mux_o_160: std_logic;
    signal mux_o_161: std_logic;
    signal mux_o_162: std_logic;
    signal mux_o_163: std_logic;
    signal mux_o_165: std_logic;
    signal mux_o_178: std_logic;
    signal mux_o_179: std_logic;
    signal mux_o_180: std_logic;
    signal mux_o_181: std_logic;
    signal mux_o_182: std_logic;
    signal mux_o_183: std_logic;
    signal mux_o_184: std_logic;
    signal mux_o_186: std_logic;
    signal mux_o_199: std_logic;
    signal mux_o_200: std_logic;
    signal mux_o_201: std_logic;
    signal mux_o_202: std_logic;
    signal mux_o_203: std_logic;
    signal mux_o_204: std_logic;
    signal mux_o_205: std_logic;
    signal mux_o_207: std_logic;
    signal mux_o_220: std_logic;
    signal mux_o_221: std_logic;
    signal mux_o_222: std_logic;
    signal mux_o_223: std_logic;
    signal mux_o_224: std_logic;
    signal mux_o_225: std_logic;
    signal mux_o_226: std_logic;
    signal mux_o_228: std_logic;
    signal mux_o_241: std_logic;
    signal mux_o_242: std_logic;
    signal mux_o_243: std_logic;
    signal mux_o_244: std_logic;
    signal mux_o_245: std_logic;
    signal mux_o_246: std_logic;
    signal mux_o_247: std_logic;
    signal mux_o_249: std_logic;
    signal mux_o_262: std_logic;
    signal mux_o_263: std_logic;
    signal mux_o_264: std_logic;
    signal mux_o_265: std_logic;
    signal mux_o_266: std_logic;
    signal mux_o_267: std_logic;
    signal mux_o_268: std_logic;
    signal mux_o_270: std_logic;
    signal mux_o_283: std_logic;
    signal mux_o_284: std_logic;
    signal mux_o_285: std_logic;
    signal mux_o_286: std_logic;
    signal mux_o_287: std_logic;
    signal mux_o_288: std_logic;
    signal mux_o_289: std_logic;
    signal mux_o_291: std_logic;
    signal mux_o_304: std_logic;
    signal mux_o_305: std_logic;
    signal mux_o_306: std_logic;
    signal mux_o_307: std_logic;
    signal mux_o_308: std_logic;
    signal mux_o_309: std_logic;
    signal mux_o_310: std_logic;
    signal mux_o_312: std_logic;
    signal mux_o_325: std_logic;
    signal mux_o_326: std_logic;
    signal mux_o_327: std_logic;
    signal mux_o_328: std_logic;
    signal mux_o_329: std_logic;
    signal mux_o_330: std_logic;
    signal mux_o_331: std_logic;
    signal mux_o_333: std_logic;
    signal mux_o_346: std_logic;
    signal mux_o_347: std_logic;
    signal mux_o_348: std_logic;
    signal mux_o_349: std_logic;
    signal mux_o_350: std_logic;
    signal mux_o_351: std_logic;
    signal mux_o_352: std_logic;
    signal mux_o_354: std_logic;
    signal mux_o_367: std_logic;
    signal mux_o_368: std_logic;
    signal mux_o_369: std_logic;
    signal mux_o_370: std_logic;
    signal mux_o_371: std_logic;
    signal mux_o_372: std_logic;
    signal mux_o_373: std_logic;
    signal mux_o_375: std_logic;
    signal gw_gnd: std_logic;
    signal promx9_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_0_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_1_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_2_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_3_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_4_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_4_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_5_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_5_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_6_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_6_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_7_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_7_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_8_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_8_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_9_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_9_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_10_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_10_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_11_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_11_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_12_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_12_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_13_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_13_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_14_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_14_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_15_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_15_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_16_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_16_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_17_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_17_DO_o: std_logic_vector(35 downto 0);
    signal promx9_inst_18_AD_i: std_logic_vector(13 downto 0);
    signal promx9_inst_18_DO_o: std_logic_vector(35 downto 0);

    -- component declaration
    component LUT4
        generic (
            INIT: in bit_vector := X"0000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic
        );
    end component;

    -- component declaration
    component LUT2
        generic (
            INIT: in bit_vector := X"0"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic
        );
    end component;

    -- component declaration
    component LUT5
        generic (
            INIT: in bit_vector := X"00000000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic;
            I4: in std_logic
        );
    end component;

    --component declaration
    component pROMX9
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(35 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

    -- component declaration
    component DFFE
        port (
            Q: out std_logic;
            D: in std_logic;
            CLK: in std_logic;
            CE: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    gw_gnd <= '0';

    promx9_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_0_dout(8 downto 0) <= promx9_inst_0_DO_o(8 downto 0) ;
    promx9_inst_0_dout_w(26 downto 0) <= promx9_inst_0_DO_o(35 downto 9) ;
    promx9_inst_1_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_1_dout(8 downto 0) <= promx9_inst_1_DO_o(8 downto 0) ;
    promx9_inst_1_dout_w(26 downto 0) <= promx9_inst_1_DO_o(35 downto 9) ;
    promx9_inst_2_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_2_dout(8 downto 0) <= promx9_inst_2_DO_o(8 downto 0) ;
    promx9_inst_2_dout_w(26 downto 0) <= promx9_inst_2_DO_o(35 downto 9) ;
    promx9_inst_3_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_3_dout(8 downto 0) <= promx9_inst_3_DO_o(8 downto 0) ;
    promx9_inst_3_dout_w(26 downto 0) <= promx9_inst_3_DO_o(35 downto 9) ;
    promx9_inst_4_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_4_dout(8 downto 0) <= promx9_inst_4_DO_o(8 downto 0) ;
    promx9_inst_4_dout_w(26 downto 0) <= promx9_inst_4_DO_o(35 downto 9) ;
    promx9_inst_5_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_5_dout(8 downto 0) <= promx9_inst_5_DO_o(8 downto 0) ;
    promx9_inst_5_dout_w(26 downto 0) <= promx9_inst_5_DO_o(35 downto 9) ;
    promx9_inst_6_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_6_dout(8 downto 0) <= promx9_inst_6_DO_o(8 downto 0) ;
    promx9_inst_6_dout_w(26 downto 0) <= promx9_inst_6_DO_o(35 downto 9) ;
    promx9_inst_7_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_7_dout(8 downto 0) <= promx9_inst_7_DO_o(8 downto 0) ;
    promx9_inst_7_dout_w(26 downto 0) <= promx9_inst_7_DO_o(35 downto 9) ;
    promx9_inst_8_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_8_dout(17 downto 9) <= promx9_inst_8_DO_o(8 downto 0) ;
    promx9_inst_8_dout_w(26 downto 0) <= promx9_inst_8_DO_o(35 downto 9) ;
    promx9_inst_9_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_9_dout(17 downto 9) <= promx9_inst_9_DO_o(8 downto 0) ;
    promx9_inst_9_dout_w(26 downto 0) <= promx9_inst_9_DO_o(35 downto 9) ;
    promx9_inst_10_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_10_dout(17 downto 9) <= promx9_inst_10_DO_o(8 downto 0) ;
    promx9_inst_10_dout_w(26 downto 0) <= promx9_inst_10_DO_o(35 downto 9) ;
    promx9_inst_11_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_11_dout(17 downto 9) <= promx9_inst_11_DO_o(8 downto 0) ;
    promx9_inst_11_dout_w(26 downto 0) <= promx9_inst_11_DO_o(35 downto 9) ;
    promx9_inst_12_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_12_dout(17 downto 9) <= promx9_inst_12_DO_o(8 downto 0) ;
    promx9_inst_12_dout_w(26 downto 0) <= promx9_inst_12_DO_o(35 downto 9) ;
    promx9_inst_13_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_13_dout(17 downto 9) <= promx9_inst_13_DO_o(8 downto 0) ;
    promx9_inst_13_dout_w(26 downto 0) <= promx9_inst_13_DO_o(35 downto 9) ;
    promx9_inst_14_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_14_dout(17 downto 9) <= promx9_inst_14_DO_o(8 downto 0) ;
    promx9_inst_14_dout_w(26 downto 0) <= promx9_inst_14_DO_o(35 downto 9) ;
    promx9_inst_15_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_15_dout(17 downto 9) <= promx9_inst_15_DO_o(8 downto 0) ;
    promx9_inst_15_dout_w(26 downto 0) <= promx9_inst_15_DO_o(35 downto 9) ;
    promx9_inst_16_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_16_dout(8 downto 0) <= promx9_inst_16_DO_o(8 downto 0) ;
    promx9_inst_16_dout_w(26 downto 0) <= promx9_inst_16_DO_o(35 downto 9) ;
    promx9_inst_17_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_17_dout(17 downto 9) <= promx9_inst_17_DO_o(8 downto 0) ;
    promx9_inst_17_dout_w(26 downto 0) <= promx9_inst_17_DO_o(35 downto 9) ;
    promx9_inst_18_AD_i <= ad(9 downto 0) & gw_gnd & gw_gnd & gw_gnd & gw_gnd;
    promx9_inst_18_dout(17 downto 0) <= promx9_inst_18_DO_o(17 downto 0) ;
    promx9_inst_18_dout_w(17 downto 0) <= promx9_inst_18_DO_o(35 downto 18) ;
    lut_inst_0 : LUT4
        generic map (
            INIT => X"0001"
        )
        port map (
            F => lut_f_0,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_1 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_1,
            I0 => ce,
            I1 => lut_f_0
        );

    lut_inst_2 : LUT4
        generic map (
            INIT => X"0002"
        )
        port map (
            F => lut_f_2,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_3 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_3,
            I0 => ce,
            I1 => lut_f_2
        );

    lut_inst_4 : LUT4
        generic map (
            INIT => X"0004"
        )
        port map (
            F => lut_f_4,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_5 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_5,
            I0 => ce,
            I1 => lut_f_4
        );

    lut_inst_6 : LUT4
        generic map (
            INIT => X"0008"
        )
        port map (
            F => lut_f_6,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_7 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_7,
            I0 => ce,
            I1 => lut_f_6
        );

    lut_inst_8 : LUT4
        generic map (
            INIT => X"0010"
        )
        port map (
            F => lut_f_8,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_9 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_9,
            I0 => ce,
            I1 => lut_f_8
        );

    lut_inst_10 : LUT4
        generic map (
            INIT => X"0020"
        )
        port map (
            F => lut_f_10,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_11 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_11,
            I0 => ce,
            I1 => lut_f_10
        );

    lut_inst_12 : LUT4
        generic map (
            INIT => X"0040"
        )
        port map (
            F => lut_f_12,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_13 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_13,
            I0 => ce,
            I1 => lut_f_12
        );

    lut_inst_14 : LUT4
        generic map (
            INIT => X"0080"
        )
        port map (
            F => lut_f_14,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_15 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_15,
            I0 => ce,
            I1 => lut_f_14
        );

    lut_inst_16 : LUT4
        generic map (
            INIT => X"0100"
        )
        port map (
            F => lut_f_16,
            I0 => ad(11),
            I1 => ad(12),
            I2 => ad(13),
            I3 => ad(14)
        );

    lut_inst_17 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_17,
            I0 => ce,
            I1 => lut_f_16
        );

    lut_inst_18 : LUT5
        generic map (
            INIT => X"00040000"
        )
        port map (
            F => lut_f_18,
            I0 => ad(10),
            I1 => ad(11),
            I2 => ad(12),
            I3 => ad(13),
            I4 => ad(14)
        );

    lut_inst_19 : LUT2
        generic map (
            INIT => X"8"
        )
        port map (
            F => lut_f_19,
            I0 => ce,
            I1 => lut_f_18
        );

    promx9_inst_0: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000C36334DB71D6DC75B71D6DC75368C633198C8C",
            INIT_RAM_01 => X"000000000000000000458000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"8EC75A68C4631918D3000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000004622C0000A534D36D300001168C6DC763B1D8ED823B1D",
            INIT_RAM_05 => X"00000000000000000000000000000000008B000000000000000000000000000000000000",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"8EC763B608EC763B608EC758CC6632322960000000000000000000000000000000000000",
            INIT_RAM_08 => X"00528000000000000000000000000000000000001A8D40000295148EC763AC361A32289B",
            INIT_RAM_09 => X"000000000000000000000000000000000000000000000000000113000000000000000000",
            INIT_RAM_0A => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"8ED82288B45B6E3B608EC763B1D8EC763B1D8EA318D4B69A6E3B1D000000000000000000",
            INIT_RAM_0C => X"000000000000000000A500000000000000000000000000000000000046A940061C523B60",
            INIT_RAM_0D => X"000000000000000000000000000000000000000000000000000000000000000000022600",
            INIT_RAM_0E => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"8E528008CB0476C0DC6E475A6C68A4763B1D8ED823B1D8EC75B9606DA3118D58EC763B13",
            INIT_RAM_10 => X"00000000000001160000000000000000014AA50000000000000000000000000000000000",
            INIT_RAM_11 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"4623228DB8ED822689000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"00318000000000011A00001A71D8ED81B89BB0476969BB04763B1D8EC763B1D8EC76C11D",
            INIT_RAM_14 => X"000000000000000000000000000000011600000000000000000112630000000000000000",
            INIT_RAM_15 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"8EC763B1DB04763B1D464523B248EC4D1383000000000000000000000000000000000000",
            INIT_RAM_17 => X"45800000000000000045B280000A50023800004323B1D8EA6DC11D8EE5A3B1D8EC763B1D",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000044C0000000000000000022600",
            INIT_RAM_19 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"8EC75B91D8EC763B1DB04763B1D8EC763B146DC75D52289E0F0783000000000000000000",
            INIT_RAM_1B => X"0000000000022C008B0000000000000000004622C00000046800C600582C0DC4EA763B60",
            INIT_RAM_1C => X"000000000000000000000000000000000000000000000000000000000000000004500000",
            INIT_RAM_1D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"69C75B8E04ED82C11D8EB71371D8EC763B608EC763B1D8EC763B148E9AA491DE560F0783",
            INIT_RAM_1F => X"000000000003280000000000000A5528008B0000000000000000D44580000004A31A94C6",
            INIT_RAM_20 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"351A9B88AC1E0F0644000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"6300000C66A466948CB0475B89DB0371B91D6E382C11DB04763B1D8EB723B1DB0476C0DC",
            INIT_RAM_23 => X"0000000000000000000000000008A5280000000000000A500000CB0000000006180118D4",
            INIT_RAM_24 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"71D823B1D8EC763BA9D4EA62844C1E0F068A000000000000000000000000000000000000",
            INIT_RAM_26 => X"00000000061801A68CA580000946209627148ED813AE06E5823B22702763B1D8EC76C11D",
            INIT_RAM_27 => X"00000000000000000000000000000000000000000000089800000000000008B000022600",
            INIT_RAM_28 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"4ED823B608EC763B22B44763B1D8EC76D06A354891383C1E0F06DC000000000000000000",
            INIT_RAM_2A => X"0000294000000196000000000006134D94C462001A6C2466C1951D4D955C0DC8EC7536E0",
            INIT_RAM_2B => X"000000000000000000000000000000000000000000000000000000000000000898000000",
            INIT_RAM_2C => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"4D955C09B8EA6DC0E04ED823B1D8EC76456F8EC763B1D8EB8CD46A353730783C1E0D1560",
            INIT_RAM_2E => X"0000000008980000000052A954A00001A800000000000A526E96C261A3196C28CAB226A2",
            INIT_RAM_2F => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"3522F0783C1E0DB91D000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0034D84C4D82B228554EA75C11D6E275C49D703723B1D8EC74D5248EC763B1D8E9AB526A",
            INIT_RAM_32 => X"00000000000000000000000000089800000000448008B0022E94006180000C465B2D88C2",
            INIT_RAM_33 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"8EC763B1DB41A8D46A529130783C1A25B8DC000000000000000000000000000000000000",
            INIT_RAM_35 => X"6180000C2EB30E954A6AB1185197A271B8DC4EB82C11D70383529D70476C11D8E9A8D51D",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000C5650000000A5000008C0035000C4",
            INIT_RAM_37 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"705823B1D921A94B1D8EC763ADC351A8D46A52E0F0783C1A2A3A89000000000000000000",
            INIT_RAM_39 => X"45800008B0032D86C40000188CB4A51226C40AB0984EA7A38E249D70381B9604EB814AE2",
            INIT_RAM_3A => X"000000000000000000000000000000000000000000000000000000000000113A50000000",
            INIT_RAM_3B => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"4EB81B9E84EA75C5A96E4763ADC351A9C71D6E476C124D49A8D46A2AE0F0783223739444",
            INIT_RAM_3D => X"00000011300000011200001A8000035688C30030D844B4631244CB6251227B075C68AAE0",
            INIT_RAM_3E => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"EBE0F07832222B06C5000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => promx9_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => promx9_inst_0_AD_i
        );

    promx9_inst_1: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"61312C6F4ADF5DC0E070275B9A94EB81C46A6E4763A6A351AA3B1DB04763A6A351A8D46A",
            INIT_RAM_01 => X"0000000000000000000000000D300000010C00001960045B2D840000309969365B4E3313",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"8ED82486A351A8D46A7160F0783C1E0C8944000000000000000000000000000000000000",
            INIT_RAM_04 => X"6230918DB6158EB6C26136D58AA4DB71C0E04EB813B2D6E581C12D6E476446A352963B1D",
            INIT_RAM_05 => X"00000000000000000000000000000000000000000011900002950C0000118C385B098400",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"6DC74D46AD4C923B1DB065F526A351AB526A64E0F0783C1E0E8944000000000000000000",
            INIT_RAM_08 => X"0000196C385B0988C36131136DB43271A6C2A5894E8A44DC993AE04EA753B7070295C570",
            INIT_RAM_09 => X"0000000000000000000000000000000000000000000000000000000000000D3000029400",
            INIT_RAM_0A => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"703813A72701A9C472CBB8F526A3538A3B1DB0288D46A351A8D46A2AE0F0783C1B168944",
            INIT_RAM_0C => X"0000001190000226000030D960065B0984C26132D38CB89B8D96C291095C71C93389C09D",
            INIT_RAM_0D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"64E0F078344D128944000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"B1CAAC8E371B81C0E070381C072715BDC4726D9AB526A354763B228EA94D46AD49A8D46A",
            INIT_RAM_10 => X"0000000000000000000000000D300002180061B0996C365B0984C26125138CB6DD6D16D3",
            INIT_RAM_11 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"8E9A8D46A351A8D46A44E0F0644A25128944000000000000000000000000000000000000",
            INIT_RAM_13 => X"62469C6C44E59227637529156EB933813AE04EB814A72715C1C6726E1A8D46AD4C763B24",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000001190030E24006230996C465B098544",
            INIT_RAM_15 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"911AB526AD4B6ED124719A8D46A351AB526AC1E0C8944A25128844000000000000000000",
            INIT_RAM_17 => X"61309974A65B0984C269D6EB6D371BAAC62552469D4B24EB81C0E07038B5272711CAD170",
            INIT_RAM_18 => X"0000000000000000000000000000000000000000000000000000000000000D30030E18C3",
            INIT_RAM_19 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"96B70D57071DC25AABD49AB526A92370D49B356A4D46A351A8D5A9C1E0D8B44A25128844",
            INIT_RAM_1B => X"000000114A531224C46130996CBA23110D4B69B4DC713ADD8EC6EA522AE70EBB0581C09D",
            INIT_RAM_1C => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"C1B168944A25118B44000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"8D4E2712693581C0A5D4A76E02C96CB65A6A351A8D52D921AADF24351A8D46A351A8D4E2",
            INIT_RAM_1F => X"00000000000000000000001894A89B1219446130996CB6134E954B45B8D3914B258C4AA4",
            INIT_RAM_20 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"351A8D46A351A8D4C944C2A8944A25128944000000000000000000000000000000000000",
            INIT_RAM_22 => X"4DD9138DB9A58D58A455BD1E960513813B7052B88E570B85C2E12D351A8D46AD49AA5BA9",
            INIT_RAM_23 => X"00000000000000000000000000000000000000001840069B0A24C26130918CB6248984D3",
            INIT_RAM_24 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"351AA5B2D351A8D46A351A8D46A351A8D489A8C2A8944A25128944000000000000000000",
            INIT_RAM_26 => X"61309968C8636D855B69B4EC75B753D1571A7A4E256EB933814A72716A65B70755C2E06A",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000030D840069B0A9744",
            INIT_RAM_28 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"6E4B6E07291DC0E5A9356A4E46AD49C8D46A969A8D46A356A5C70A71D128944A25128944",
            INIT_RAM_2A => X"00312880069B0A96C26130996CB8CC4D1894ADD6C4ADC9C4E2352A9C4E155704ED82E072",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000C3000018800",
            INIT_RAM_2C => X"71D128944A25128844000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"9C4E154EB70296E072B01CA5A6AB45C2E1A9354B6E06A355C3532D351A8D46AD49ABAEE3",
            INIT_RAM_2E => X"0000186D5000010C000031184C389B0A94C26130996CBB1C4E32946DB8D38EB9C3B136F4",
            INIT_RAM_2F => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"351A8D5A9351A9C66A855468944A25128903000000000000000000000000000000000000",
            INIT_RAM_31 => X"68B8D39349C591B9387A4E1E9224EDC2E0ABB45C0E49B395C25A6A355C2E1A996CB75370",
            INIT_RAM_32 => X"0000000000000000000000116E30000184C30030984C489B0B2CC26130996CBB1A31B69C",
            INIT_RAM_33 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"96DC25A6AB81AA5B70D49A8D46A351AB52E3A22528944A21120703000000000000000000",
            INIT_RAM_35 => X"A251196D34E44EC6DAADA71B8F47A29156F49C4E164E052DC1D52DB85C0D560394B4D46A",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000119A96180288C30051184C20032E94C2",
            INIT_RAM_37 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"B85C14AA5B81C8D46AB85C2DF70166A65B2DD49A8D46A351A8D5514A38E8944A240E0703",
            INIT_RAM_39 => X"0030984C20036E954A6130996D34E465389CADD8EB6F45526DE9389C4E154E0B79CA4970",
            INIT_RAM_3A => X"00000000000000000000000000000000000000000000000000000062D29966ACB80312C2",
            INIT_RAM_3B => X"B8252894481C0E0703000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"9C4E144E2B84B5C570B85C1B82CB81A8D472B84B65B70969AAE12D351A8D5A9351A9C70A",
            INIT_RAM_3D => X"62B29986A7152F2F856230A88C26234D854A61309971A4E58DC694ADA72B73871B8E7138",
            INIT_RAM_3E => X"00000000000000000000000000000000000000000000000000000000000000000001A200",
            INIT_RAM_3F => X"D49A8D4723538EA2E396D10890381C0E0703000000000000000000000000000000000000"
        )
        port map (
            DO => promx9_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => promx9_inst_1_AD_i
        );

    promx9_inst_2: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"ADA71C7384DAA9E8F49C3D244EAB8295D57096EA5C570396A6E170B84B6E12D355C2E1A9",
            INIT_RAM_01 => X"6500000000022D8A9242B2D0A6A52B7296556151288C26144D894B613090C9C4E58EB694",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"B85C2E12D96DC2E06A355C0E46A3575E5B7085112070381C0E0703000000000000000000",
            INIT_RAM_04 => X"61512969C4E58DC69369A7156AC722B271389C2CA44723965EE17039277532DB7CB6E170",
            INIT_RAM_05 => X"00000000000000014A62B2994CA0033196CB663460AE335382269DA261712C2A2312294A",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"D4B725B7096DC2E170B85C2E12DB85C0D46A161C8D46A71B8EE0E381C0E070381C0E0703",
            INIT_RAM_08 => X"4EB09B8C261309A74A6130A271A71A71C6D36989669348D4E271389C2A8D02C9226EE170",
            INIT_RAM_09 => X"00000000000000000000000000000002940065248009262B2996CB65B2D491C35295C09D",
            INIT_RAM_0A => X"81C0E070381C0E0684000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"9C4AEE4EB71296E07271380E570B85C2E170B85C25B2D96CB6DF70B81A8D4E3165C1B703",
            INIT_RAM_0C => X"68A6E35A5351A9C09D702753AC261511A8C2A530A329469A4AB69469A71D91A55BD27138",
            INIT_RAM_0D => X"000000000000000000000000000000000000000021800003158A856632DA28568D2996CB",
            INIT_RAM_0E => X"B7B8CD57096A52150681C0E07444240D1786000000000000000000000000000000000000",
            INIT_RAM_0F => X"69B71E8D9D84E271389C3B1D7704E9AA5A6A4EA965B70B85C2E170B85C25B7096DC25B70",
            INIT_RAM_10 => X"42C2D96D165B2D96CB65E9546AB356A4D49D4EA753A8B65B0A94CBAAD111893AB4292556",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000022C01146500116D1",
            INIT_RAM_12 => X"96CB6E170B85C2E12DD4CB6E0AB65A298AC581C1A870681B2E0A4B000000000000000000",
            INIT_RAM_13 => X"6130994CA49A4812D349A5159569C2B1E938563AE49A96E4B4E4E24E9A9D570B84B6E170",
            INIT_RAM_14 => X"69801A74A6A31A94858541686C665B2D96CB65A48E4AAB86A4D4E24EB813B1242B0984DB",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000C40000000000000000000000000D3",
            INIT_RAM_16 => X"6E5A0E570B85C2E170B85C2E170B85C25A6AB85C0D5124531289038350D8884653188F03",
            INIT_RAM_17 => X"B03813AD365A2D0AD4A530891436232C049365329D493562B270AC6D275C6E2701C8D49D",
            INIT_RAM_18 => X"0000000000031694006DB6E968C4DD2A958665C18130A6332D96CB65A4F4B2DB85C0D46A",
            INIT_RAM_19 => X"A1D120D0565B2A07030000000000000000000000000000000000006180000CB000000000",
            INIT_RAM_1A => X"4EB80D49D529C9C4E071296E170B85C2E170B85C2E170B85C25B70166A5148A628098B06",
            INIT_RAM_1B => X"632634A2C719CA5A6A35274AB1362B2C89444DB2E160245A4C040385C174698D1AB1591A",
            INIT_RAM_1C => X"0052C0185A500000000000000000030E28DB464762960CB34E949265828040204B1996CB",
            INIT_RAM_1D => X"5295614C501D1109440111D94CB82A2A07030000000000000000000000000000000000C3",
            INIT_RAM_1E => X"01B1930D168F69A3604EA77D09D529A93A9DB03AAE12D968B2E170B82AEE17096CB6E170",
            INIT_RAM_1F => X"8500805446200D0AC66561B4B2DB826EE06A35388ABD76591289C8C33149003014280402",
            INIT_RAM_20 => X"00000000000000008C0032C0185428000000000000000A552987608ED82C1608EB699786",
            INIT_RAM_21 => X"B84925B70B85C2E0A56E12A0D440191D8A02A222D8CCB62C0E0703000000000000000000",
            INIT_RAM_22 => X"65D11960305008060301D0C12D165B45A69D4EA75C49DB8371C0E0701CAE170B81AADE2C",
            INIT_RAM_23 => X"B03932CDBB04750B058500C0402623120ECB6532C90F23428AE170D49A9361565B16884A",
            INIT_RAM_24 => X"0000000000000000000000000000000000C6A2625968544B10000000000008B004522996",
            INIT_RAM_25 => X"711CA5A72B7A6CE570715C2E170B85C1D49D64C0D8802A2418040245C1596CB4240E0703",
            INIT_RAM_26 => X"969A946CBA25128944A21121544013640447A211C12CB65B2DA69B4EB813A9DD4B81C0E0",
            INIT_RAM_27 => X"0032C00008A00137608EA88E4DBCE581AA93850080402A231488446211094D53438D3672",
            INIT_RAM_28 => X"82B2D970781C0D08C500000000000000000000000000000000014B42A17068562A140000",
            INIT_RAM_29 => X"703813AE2B03813AE0D4DC2E1A96E1AA5A6A925C2E02C96CB53A9D85212860223B100544",
            INIT_RAM_2A => X"6251288CB7567338A2391AA468BA241E8944A251188C4A259407066240D0A928D32D969B",
            INIT_RAM_2B => X"A5224898364E0D88000052988004634D191DB0476483451673C0D445D10040A8311D8A44",
            INIT_RAM_2C => X"81D10040262008054465B2D968442315888B0000000000000000000000000000000000CB",
            INIT_RAM_2D => X"23C0C069BB937196D3B4581C4DC71275C09D355C1C49D6E1CA5ADC968B2E02C51B713B12",
            INIT_RAM_2E => X"6A22C96478340E0684832108913CE38F3955750B14744623158B44A211188D9A25960C47",
            INIT_RAM_2F => X"0000000000000000C344E1512C562B1488C30031114C6AAC75B71D8EC763AABB858338DB",
            INIT_RAM_30 => X"96DC25B5671A753B0A81808040201808060965B2E890AA202A16C6000000000000000000",
            INIT_RAM_31 => X"A236EAC7B792AFA90A81C0E0D261A24D311A753894AA571389C09D39389C09D354B6C0E2",
            INIT_RAM_32 => X"B05823B1D395C1B7E0CE32E0D038540E07034240E06CBCE673C16089392160A65E118AC5",
            INIT_RAM_33 => X"000000000000000000000000000000000000C2A17094422510888A0030CAA8B8A4523B1D",
            INIT_RAM_34 => X"71381C0E2B85813B6F96CB5550B6E274AB036200804020180804C665B2D174301C1596CB",
            INIT_RAM_35 => X"4E32C060262E0D8A4AA25126F791D8EE4CDA81C0E0D261A291491C55C92DEEA7138B529D",
            INIT_RAM_36 => X"450011513E54763B1D8EC75C6DB724B76755CE557A70A81C0E070381C0E07C98A26F399C",
            INIT_RAM_37 => X"6350C04096332D9706000000000000000000000000000000000000A560C88C5A25121583",
            INIT_RAM_38 => X"555BD5770755A14A9D703813B6F6E275C570390B288CB4EB809503010080402010090ACB",
            INIT_RAM_39 => X"8542A070AEA35339E06AC1A8707629119294A212996A355A4D3172EA40E06DA553C98CDC",
            INIT_RAM_3A => X"61A258AC5A251288C5C1A2B959789E5EC11D8ED8144AB6DDC2E068CE781970381C0E070A",
            INIT_RAM_3B => X"0100804020180C12C68500804C665B2C128B000000000000000000458000000000000000",
            INIT_RAM_3C => X"9342A06DA1A595A292791CAE17055DC1B9A96E38AC09D4EA765B701642C07127027614C5",
            INIT_RAM_3D => X"CE782290A8575196CB63121170A81C29A79C8A42807C8429118AE34A2525A2C69B691764",
            INIT_RAM_3E => X"A531400000000186CB002150AC9A2512890AC1F2912558EB723B1D8EC75C8E3B7B92E072",
            INIT_RAM_3F => X"45809969D7044A07440100804020100D8D430100C12CB65B181402000000000000000000"
        )
        port map (
            DO => promx9_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_5,
            RESET => reset,
            AD => promx9_inst_2_AD_i
        );

    promx9_inst_3: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"3938C587255C1E06CB45B2D38EB8D24924EB75DC2E12DB838EDF68D4B89C09D4EA96E02C",
            INIT_RAM_01 => X"B04763AAB55DC2E1707278225D424000014A665298AC68540C975969C288EC544A168951",
            INIT_RAM_02 => X"00000000000000000062B280000000000085A23098AC562D1289C8A8E12268A8EC763B1D",
            INIT_RAM_03 => X"B4275C0E04EDC3AECB0100A269D4E9298A020180804020100A86020121596CB630240402",
            INIT_RAM_04 => X"45C0C8F84A232E0ECB519C8E4348D36E069471581A6000052A687B793AEE52DB81CAD0E3",
            INIT_RAM_05 => X"65D44AB136E4763B1D8EC7544E3164B65B7039557388C0032D24CB65B45974A61C2A14D5",
            INIT_RAM_06 => X"A1B199609010080402000000000000000000A5528000000529874A2262688C5A2512884A",
            INIT_RAM_07 => X"593CCE8F296DC2E06A6E3813AE07144D26030122DB89D2AA2A89060180804020100C0402",
            INIT_RAM_08 => X"62B1596D142B2E070725C290A89431210ACA6528CE4341A0D1B7C84EA6E3B4B005C9E67B",
            INIT_RAM_09 => X"64E118B4462D12894489C52271D6E5823B1D8ED81C6EA91DC2E17096C72254A68B2E9485",
            INIT_RAM_0A => X"A2008040201008040204B2D0A03010080647000000000000000000A541400000000234C3",
            INIT_RAM_0B => X"4EA75B74B8E5E476B43D9EE70B2795C8E4EA353893A9D89A2E8603A244D369D8531516CB",
            INIT_RAM_0C => X"B81C8000062D2A954A42A150B05688021506852290AC4A521596938E1C868341A1C8690A",
            INIT_RAM_0D => X"65B2C000000001C6CBC2B258B4462D128944A8C7628DC8EC763ADB8EC763AE4B85C2E170",
            INIT_RAM_0E => X"4644DA6DC4542E26C40180804020100805436302404020100A888A000000000000000000",
            INIT_RAM_0F => X"D9DC068341A0D0688A2AE5800DA9B8ED68353D9ECF738763ACE52D55C9226CBA20080402",
            INIT_RAM_10 => X"B036DC6DB55DC2E170B85C1AB4A0032A954AA53290B4A65D28970381F228800A5347B51A",
            INIT_RAM_11 => X"00000000000000000068B2C00C50030DD868C2B2488CB225128944A244DB9608EC75C722",
            INIT_RAM_12 => X"6632C120201808050B65A2E24CB45C4E26020100804020100806096302404020100896E3",
            INIT_RAM_13 => X"8521400CA65B2D8CA3969C868341A0D068D571625AA723D8EC767BBCAE8F67B7A5E6E5A5",
            INIT_RAM_14 => X"A2429B71DB0475B6EA6DB8DC6EA8EDC2E170B85C15400A53150ACA00215A2CB65D299703",
            INIT_RAM_15 => X"0100804030122DC6F40000000000000000CA65B2D1600A5001D8BA453158AC565D119744",
            INIT_RAM_16 => X"759ECF6B81B2CB4BA58D32D0B0A0100806CB85B2CABD68995616020100804020100E86C6",
            INIT_RAM_17 => X"A532D96CB65D29970345D28014A65B2D97A5B84B469371A4DC69134EE5DB4F21D9EC7665",
            INIT_RAM_18 => X"95612884AA512996CBA2512271D8EC76C0E355C75D52355B92E12D96CB4E4E38A5280000",
            INIT_RAM_19 => X"0480804020100E0A090180C04020538DE93800000000000000014A65C1694C562B14F67B",
            INIT_RAM_1A => X"A5B71C9B3BC8EC767B8E2ACF67B3DBD3B4926332D1543A180804030526DC48B2AA300456",
            INIT_RAM_1B => X"B82AF66F28A45294D568B2D96CBA552996CB893AE94CB65B455570968D068F29BAD2F2EB",
            INIT_RAM_1C => X"65D2996CA63329747B3DC7115444A32C94CBA8D1095978EC75C6DB55BA936AB755C2E170",
            INIT_RAM_1D => X"89B8227D74A00E14340100804020100A86020180C0603B23D270360000000000000000CB",
            INIT_RAM_1E => X"51F5EE4B479DE6707B75D2E46F2BC9EC767B9BB6ACAAA3D9EDA2D16332C1305048080403",
            INIT_RAM_1F => X"8EDBE5AEAB85BEE170B81C9A665D2C51394A6E32E954AA552801141B34D96CB65AAAE0E3",
            INIT_RAM_20 => X"0000000000000000CB65A1596CA62A4974AA3DAEA39448556626CBA542A88CB8EC763A72",
            INIT_RAM_21 => X"04A2915430100806CB4532D16CB45D0D56560100804020100A89440180805DA9C4E158DC",
            INIT_RAM_22 => X"6DB4DA2CB8D28EA3444A156F2BA3DAE8F67B3DB4DD572BC8EEF23BB932E14E4343B196C6",
            INIT_RAM_23 => X"6D34EA2448A4763AE4392AEE07296DC2E0AB164B4D1194E27350DB00316954A65315C6EC",
            INIT_RAM_24 => X"0180C2AF47A3AD3603000000000000018AD165A1412CC42A4975A39C271D71C65A533912",
            INIT_RAM_25 => X"3D9A118D9340D7B4D16300C04020100804CB45C2D969B04D94F6090180C0602A23111602",
            INIT_RAM_26 => X"5936E94CA89C893919B1A49A2CB5232E8844A2371D4BA3DAC8F7383DB6CD0721D8ECF63B",
            INIT_RAM_27 => X"1468DB4E334546AB5589B6EAB12A8C52C0DB96DC25B70B85C25B2D6DE974B19594E1E938",
            INIT_RAM_28 => X"0100A888B4580804020144D58EC5244C040200000000000001949204D2996CBA532DE7A3",
            INIT_RAM_29 => X"5D528E5793D8ECF722BC9EE39C9951EF47DA65A280403015108EC401C2D3656B29EDE402",
            INIT_RAM_2A => X"3946538F49C4E1E9387A4E1E8B2756A2C763B1A49A2CB6532E88C5A22753AEB3DD8CF6EC",
            INIT_RAM_2B => X"4541514CB68D2BB5DA688A1A76032B56279CCE355B7554A2532CEA8EBAAE170B82ACE472",
            INIT_RAM_2C => X"A1D96CB2B1D8EC140201B11C8030100C040201E8E54E38500C0403005280000000010ACB",
            INIT_RAM_2D => X"852753ADC9A09564EA7647058F2BC8ED692A719EECBD625CA954CB65826874423B100403",
            INIT_RAM_2E => X"721CA5B70B83AE24E38CEA256B2756A1D4EA750944A2512896C625B1B45A2CC65D1288C9",
            INIT_RAM_2F => X"0044C0000003299609048250ACB6332D961568F69A2E39265A289BCE6733860CE5553714",
            INIT_RAM_30 => X"82C2D170BA251288D91A2ADE47B3DD95888B62594AC030502A888B4DBAF4713018080402",
            INIT_RAM_31 => X"B1D8245136591215122AA75C16091095D963B1A8D462C794DCF6E3B22D0AC84424A86428",
            INIT_RAM_32 => X"B0673C19CCE7833996CE554D0EBD9DC9692B7A3D165128CA704B63B18944A2512D8C4B63",
            INIT_RAM_33 => X"5668C12020100804090032A291200345968A63215140904B2D8CD104F6996DA355BF2C9B",
            INIT_RAM_34 => X"959EEF2C581CAAC89885B29168B6CC9A56341A0D256E47222C0402B2D96870B6CA2D16E3",
            INIT_RAM_35 => X"B1D8EC763B1896C763B1C8941602AD1288552AA75C16012D8C4B63D1A2D46A3D9BC87770",
            INIT_RAM_36 => X"04B2D96D3F46A6DF96CE673C060F078339E0F0283C0A0D83D1E8B2594662512892735025",
            INIT_RAM_37 => X"7222DB326A2027B4AC0A80C04030100812AC6AA6DC6D469B2C128A04C281343453199609",
            INIT_RAM_38 => X"ED009470B390B1E5374E3C8772681B50D09845A4D269C934AE4D2B95CAEE4344980A8965",
            INIT_RAM_39 => X"8944A25128CA72C76312D8C4A2512D8C4A2512C89C71D4DC2A149D2AB813B60B1D8DD4EA",
            INIT_RAM_3A => X"A180D8C0342A15968A4532D96D1911AB526A6DE73C19CCE6733860304AF51B07A4E35119",
            INIT_RAM_3B => X"95CAE56E449B65C8E42B5C8F6560576B46090100804020102B47A369B2DD5138A34594C6",
            INIT_RAM_3C => X"4EA76C160D43A9D4F4D180A160A45A8E3472B938E6EEB6D40D36CB85B2D96CB8A42DA72B",
            INIT_RAM_3D => X"CE78256B29C4E3611289529888C89466C76312896C763B1896C763B1A71B7606E3251255",
            INIT_RAM_3E => X"69C5164D38CB2D96CA04A150A0204D0D968542B2D96CB8EEA4D56FB438F399CF0670C19C",
            INIT_RAM_3F => X"4A26D369B723C9552BB95CA56561A0D0D765BC8EECA0945054060201808040204F6958E4"
        )
        port map (
            DO => promx9_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_7,
            RESET => reset,
            AD => promx9_inst_3_AD_i
        );

    promx9_inst_4: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"D438EC1608EA6FAE9D7027644E3B1ACA70EAD180805440124D26AA55BAEE4344E40E06DB",
            INIT_RAM_01 => X"B065B39E0F078339E030672B3198CA8232C365D47AF128CD8E45A8B1896C62512D8C4B63",
            INIT_RAM_02 => X"010280609ED2B064E38CC51D5638A32D9706A180E86850100D8D4342B2D96D16D38F52DC",
            INIT_RAM_03 => X"3946859707592E070A4A5823B1D8EE965579BC8ECF63B1DBC8F63B1D9EE870A048080602",
            INIT_RAM_04 => X"B1D8EC625B1D8C4B22B04763ADC8EB71B89D6E48AC060B1BAA70F47A024040201D11391A",
            INIT_RAM_05 => X"4282596926D476486A351AAD0DBCE673C19CCE7833959894319751A21118C8C6DA51A69C",
            INIT_RAM_06 => X"1D82404038515814022B02812157A4E1E8F312C66C6F48CB2D96CA83808070A010091402",
            INIT_RAM_07 => X"557680402018091770B846B4B70D9D5A0703854523B1D8ED834A74BC8EC763B1D8EC763B",
            INIT_RAM_08 => X"8532F911389D2A3225B18953963B189645608EC763B1D8ED823A9BB0181C6E3B1BAB61A8",
            INIT_RAM_09 => X"83D12888501008068501A15A2D16A582D1A9351A8D56FB4477399CAA982AB12A5B2C8944",
            INIT_RAM_0A => X"BC9EC763B1D8EC767B6C8268656959A004566C827B4F49C2B168F359465A6F4B1B4D96CB",
            INIT_RAM_0B => X"CB58141225528351596E76814020100E1756B80B1A370B83AE150381B2E29608EB91E537",
            INIT_RAM_0C => X"75556188B64D128944A24290A8AA5C484B63B1C4AC76371D8EC11DB04763A9BCB3AE3B1D",
            INIT_RAM_0D => X"7A58E28EA5945196CC65B14054401008040201A15A2D16D476486A351A8D4A2755BEDF68",
            INIT_RAM_0E => X"81C2BAC8C8A451A71C32DE4767B1D8EC76B489B64F779B2826CA3404F6A70F4590EDD8F4",
            INIT_RAM_0F => X"8EC763AA2BCBC8F67B9BE73399CCE183C0DA698242A090100926CB55CB5462C161C9B903",
            INIT_RAM_10 => X"351A9D4EAB1C89C7228CB6D1584855119344A260D134B896A04B22894664460B036EC11D",
            INIT_RAM_11 => X"ED2B1D8B41A3ADD8AB563D139637A27197866511188020180804020100D8CD46D36DB768",
            INIT_RAM_12 => X"725C1D6A3B84B5D70381A3197D6EB34D4615795CAE572B95E6F2341A1EC776585D94690A",
            INIT_RAM_13 => X"8CA81371DB05823B1D8EC75B6683D9EC767B4DE70C1E0CE26E27558580914020100A88A3",
            INIT_RAM_14 => X"015110AD58D4763B1DD49A9D76F916A2C7636DC4C88C562A1688C5C1A26971212A722512",
            INIT_RAM_15 => X"6D391B353724AECA93522AE57A54C26E56E4B1EC3509C753D1A6CA6531588C4625100544",
            INIT_RAM_16 => X"6980C1202010080493559C8E4DB718B0588A81B2E291D0AB2D37266D369B4DA6D3524CDA",
            INIT_RAM_17 => X"2252A25228CC4A24D3865563B1D8EC763B1D8EB70D07B1D8EC76658A67339E0CE45234D4",
            INIT_RAM_18 => X"6532C88446231004C40150E16D36DD823A656DA8AE57075D8C4B636AB2C898362D110B83",
            INIT_RAM_19 => X"51CADC8E493499C92672271C8E472391272A95CAE56A455CAE57656A58C4BA84E3D2C6D1",
            INIT_RAM_1A => X"4A52E959C4DB4D94028300C04030100804028E48E5A9C6DB8C590AC326DC8158A38D36D5",
            INIT_RAM_1B => X"6DA2888C5A23159383C4C4A3312895563B968ED823B608EC763B1D8EB6CF63B1D9EDE54B",
            INIT_RAM_1C => X"E4B504A25D43A958D3653088944A211188C46251216936AB6E3AE3592AA5738592C84B63",
            INIT_RAM_1D => X"0AB8E28944DA6D36E4CB5C8F634B94AE576595CAEE53755A9068347938E547BB90D2F364",
            INIT_RAM_1E => X"8EE94763B1D9EE289465D45479C8D50E1602010080402010080402499AAE02C45B8DC6E3",
            INIT_RAM_1F => X"D83D2713875096C6DB4561089448531706858644A24CA6DD82C11D8EC7536DB8EC763B1D",
            INIT_RAM_20 => X"359EC767B1D8ED58B2EA725A7631289760D34930B0D44A251188C46251128D5B036D44E3",
            INIT_RAM_21 => X"A265F672D518B1C6E371C7154B25536DB49B51E965634BC8EC687BB95CA572B95CAE56A4",
            INIT_RAM_22 => X"6D352271D8EC763B1D8EDE4763B3DB92A2CBE451196CB2400804020100804020100C0543",
            INIT_RAM_23 => X"62312171D8ED823AB2D84E271387A096C71489A16154462911134B8943294DB6DB563ADB",
            INIT_RAM_24 => X"3D8ECF7791A1EEE52B95CADC8E4B938DD8AC6234D28CB8D58D382569B2D0B44A25128844",
            INIT_RAM_25 => X"0100806020100804850144E4472B848D56E30AA6D492A762B1D6E3D2C6A6F2B95B925772",
            INIT_RAM_26 => X"89249A6D449351954AA5529A9608EA6E3B1D8E9EC77797932C948C2240D150A855100402",
            INIT_RAM_27 => X"4E2498444A251094C52211188948EC763B2B9C4E270EA75095B4D44531689C8629119712",
            INIT_RAM_28 => X"955CAF27B1A1EEF32B72392572B1A0D0F779BC9EEF37975AAA54F2A530E17D6658563563",
            INIT_RAM_29 => X"2240E068481B2D16020100A88020100804026342DC4E4B838CD4E30AB69C6AC55CAA5434",
            INIT_RAM_2A => X"2251214C5C1A16254A68B2DA2D165B2D254AA552A291469C4D9723D2DE6E47B4A5440186",
            INIT_RAM_2B => X"0052A250C8592996154934D96CBE472288CBA242B90CB8A5823B60594E1E8F49C0964513",
            INIT_RAM_2C => X"B426CCAB29C3D1D96455DC8F67B1D9EC763B3D9EC697295AAECB65958D0D7A375DE568AC",
            INIT_RAM_2D => X"9BDCB66686580000CBEB40E064B83B519707A222F0CC401808040242C2936E3B7B8D29A9",
            INIT_RAM_2E => X"95CE2713812D8DB783E431489832252E949265B2D96CB6332E954AA534F930A65A3214CB",
            INIT_RAM_2F => X"55D925772B94A9C6AA0000000008630D184A65B29968C65B2E15C8C3317911389B72C160",
            INIT_RAM_30 => X"A1B1A34EA71DBCD4E351476C8DC563D1E8F4563AD48ABB93C956341D8EEF2B4192D0F634",
            INIT_RAM_31 => X"42B2E07034540D9694753C9E54B00000008646229155325A51B7856261B0C85620080402",
            INIT_RAM_32 => X"45B2D96CB89C76C0AA7A2CA70F4B1D8D178344E0C898342C49A34A65B2D96CBA552A94CB",
            INIT_RAM_33 => X"358C9E6B41D8EC77791D8EC7734563D2683500000000089432950C4612B92CA436258586",
            INIT_RAM_34 => X"42E1B91836280E86020102634A271EA4D4E351B8E56EB953B1E9385C2E06CEC55AAD56F2",
            INIT_RAM_35 => X"65B2D974AA552994CB45C0E070381C0F9294B82ADD4008A272C71461B2D14D4EA34DC6DA",
            INIT_RAM_36 => X"8643196CBE4B2E14CBA230A8944C2A29C6656D3B27025B1B6F0689C4A250A89A5C4994D1",
            INIT_RAM_37 => X"7A2B06CB83D9ECF6AB953CA57721A3C8F63B1DBCDE8363D9ECF67B00000000000000010C",
            INIT_RAM_38 => X"758020E8AE9D6C4B63226190B83C1B2D0A030150D96E475288D4EA722AD64F4562AD56AC",
            INIT_RAM_39 => X"8A3130B898634D96CB65C15974AA512114CB81C0E070381C2A14D3B7DBDAB1395AE8F67B",
            INIT_RAM_3A => X"0000000000000000000030E18C3A5B2D19514A129968542A15148A71BD1D56312C5226C4",
            INIT_RAM_3B => X"B83AD56F47A4E254AB55CE0F67B3D9ECF6BA5A2D0D6AB1A2AD56A471AD064355D1ECF67B",
            INIT_RAM_3C => X"355BD86259C3D1E8F49C4D00084E9B8C4A2545A270783C19128885018258D1C345A2D06A",
            INIT_RAM_3D => X"564E1593812C4D17128652D1512A534596CB65B2E954AA522A070381C0E070381A2EAD14",
            INIT_RAM_3E => X"190C8D66B951ACD6EB000000000000000000A534EC196AAC4986C34332D971365C491760",
            INIT_RAM_3F => X"01008129235289C66AB83D1D868563D1E836951AC6A7B3D9ECF67B3D8D5743279BCC6A32"
        )
        port map (
            DO => promx9_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_9,
            RESET => reset,
            AD => promx9_inst_4_AD_i
        );

    promx9_inst_5: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"81C0E070383B158B23351A800F475096C7637A4E1390725B704A9C6AE0F0783C1A1596C6",
            INIT_RAM_01 => X"8944A250C8643228AA9C4E271B012896251289452971268B2D96CB65B2E94CA4540E0703",
            INIT_RAM_02 => X"3D9ECF67B3D9ECF67B3D9EC6A7B79BB1593400000000000000000000319A6DAB04522512",
            INIT_RAM_03 => X"6A9130783225458A8A4280A8705B7BA9D56075CE1E8EC953ACF7389C3CCD72A191ECF67B",
            INIT_RAM_04 => X"65B2F0C4B81C0E070381C0F93076534DA92DD4C9294EA12D8EC76312AE174CB455904B63",
            INIT_RAM_05 => X"0000000006DA6EC11DCB44A199C86555C7387A4E1E82512D2A950C8952A24CB6632D96CB",
            INIT_RAM_06 => X"3D9EC6A32359AC6A7B3D9ECF67B3D9ECF67B3D9ECF7389C1ECF67B000000000000000000",
            INIT_RAM_07 => X"B1BD174D34524EC62565F2B0783C1A2496CB65D0C04CB8E1A944EA8A2C970F4562AD48F4",
            INIT_RAM_08 => X"8943226D342B2D96CBA5345148481C0E0703E492DA6C565351C86A3526D9425B1895E8F4",
            INIT_RAM_09 => X"00000000000000000000000014A864323ADB8A36E3B96AAC7564B2D84E1D4EA8A52A194A",
            INIT_RAM_0A => X"6E26DE8B83DCE1566B551ECF67B1AAAD56AB1A9ECF67B3D9ECF67B3D9ECF67B3D9ECF67B",
            INIT_RAM_0B => X"D4A6D9425128D9E8F4D83A8F6DB85252C69C8A11307832231514CB82A140609499A94A9B",
            INIT_RAM_0C => X"9C3D164B29136C0112A5432294A68B2D96CBA532D95C981C0E07C9AB3198A8B8E390686A",
            INIT_RAM_0D => X"3D9ECF67B3D9ECF67B0000000000000000000000000000034DB69B6DB6DB6D3B0581C6E3",
            INIT_RAM_0E => X"66318068A65B8DC6DC89A2E34EB7A2E0F734559A1E67B3D9EC6A6B559A0647B3D9ECF67B",
            INIT_RAM_0F => X"652158AF26D4B6E06AD4C52942512B8E32EA9C3D1709CEA24E289C6AE0C8983C1C2988CB",
            INIT_RAM_10 => X"8A582C1968EC76C1B07A3D1E9B07A52A954A0044A24CA65B2D974AA52160F034532DA8D3",
            INIT_RAM_11 => X"1A8C8D66B190D4F67B3D9ECF67B3D9ECF6B80000000000000000000000000000000000D3",
            INIT_RAM_12 => X"69B259383C1A26150A42B2D0A8565A6D37D745A294465594E06CB89C1A0D6321A9ECF67B",
            INIT_RAM_13 => X"65B2D15C9C334D8CC56322E349B55CB4E46A3526E29639BCDDD5387A3D0F6DBEA26E329C",
            INIT_RAM_14 => X"000000000000000000005823B1DB0475C738596A165B04E00000008944994CB65B2D9692",
            INIT_RAM_15 => X"3D9EC6A6B358D4F67B3D9EC6A32951A0D6323D9ECF67B3DAE1E8F4000000000000000000",
            INIT_RAM_16 => X"9C3D0F6CBEA346289C69D1306C9C1E0C97036632C128565B29288944B2CCAEB5A1ECF67B",
            INIT_RAM_17 => X"894320ACB65B2D96CB65F5216C562B310AC64521AE0DA1A5C2E06A3544E949C9B9D27138",
            INIT_RAM_18 => X"00000000000000000000000000000000000045C763B1D8EC7554B271DC1C6AA000000000",
            INIT_RAM_19 => X"C1F29B4ABD82E8F67B3D9ECF67B55AAC647B3D9ECF67B3D8C8646B559AD54369C3D1E8F4",
            INIT_RAM_1A => X"355A1949C9BBD271389C2E17448A9A4E33198A1298B44C1E0D970345D29970A65B1888C5",
            INIT_RAM_1B => X"71B8CCA0000000014AA5001A2CB65B2D974A4A30D8AC562B158C8AC2C72E1A5B85C2E06A",
            INIT_RAM_1C => X"762AE54A4524A86436000000000000000000000000000000000000A5C763B1D8EB6D5560",
            INIT_RAM_1D => X"85215968565B2D974464E0D14659A4AD747B3D9ECF67B3D8D6546B191ECF67B9C4E06CEC",
            INIT_RAM_1E => X"A25C0E4E4969CAE12D351A9869C554E271387A4E1C693A9B2A29148CC4D8B44223161503",
            INIT_RAM_1F => X"89E5A3ADB8EC76C160B0475A6000000000000032996CB65B458AC6630018AC545B191244",
            INIT_RAM_20 => X"954A86A7B3D9ECF67B3D9EC6A3595291389C000000000000000000000000000000000000",
            INIT_RAM_21 => X"8CB6E154462D458B0A81B31960965B28894442E0F068595CD1D5343D9ECF67B3D9ECF635",
            INIT_RAM_22 => X"003158ACB6322B07834DCB4E4A339492E06A351A9AAD3D40DA70B81B2E995D4A9829A69C",
            INIT_RAM_23 => X"0000000000000000000026E289B8A4763B1D8ED8294000000000000032D96CB49314014A",
            INIT_RAM_24 => X"762E8E9343D9ECF67B5D0C8D72A1A9ECF67B5D4D0E970B83A9C6E3000000000000000000",
            INIT_RAM_25 => X"3DBAD97D345A2E29146DB6E2744A2215890A81B2E94CB65C168944A260F078389ACA68EB",
            INIT_RAM_26 => X"62B2D96920000000000032916C442E0F078371DC0E52D35296E170353AAE000B1BCCF67B",
            INIT_RAM_27 => X"00000000000000000000000000000000000069A32188CB036EC0608EB6D1800000000000",
            INIT_RAM_28 => X"A2317078322695E6EC9A6A26972B91D174BA3DCD268AB4E4AAE57055BA8D46A351A8D46A",
            INIT_RAM_29 => X"351AAE09BA5095747B5D32BA7D301C2CCB146DD823B0AA221615068191E94CB651208944",
            INIT_RAM_2A => X"8EB6DB60000000000065B2D9600000018600005130A8A2260F068991DC2E17052A965B70",
            INIT_RAM_2B => X"75BA8D46A351A8D5A9000000000000000000000000000000000000000011955CE36EAADC",
            INIT_RAM_2C => X"81C2A950565C1C8944A251089832222AE0BA562E9D92BB93ADD5703A1D0E874B9695C6A3",
            INIT_RAM_2D => X"EBDC2E0726E388E570969AADE724652AC6E36522FA7D301C2CD119B04763B12A21298906",
            INIT_RAM_2E => X"0000116DB89566C19CB0475A60000001868A66331888C000000000631111583C1E0F0712",
            INIT_RAM_2F => X"351A8D4EA755BE46E371B8DC7A9351A8D46A000000000000000000000000000000000000",
            INIT_RAM_30 => X"4DC763B148540F930381C0D96CB82B2E8944A25128844C1A2B4AAB3DAC964BA594AEE52D",
            INIT_RAM_31 => X"45E0F0783C1913068971B8EE12D4EB80E4ABB83A8E47255B0C00CC0554FA7D30524DC8E3",
            INIT_RAM_32 => X"000000000000000000000018600A526F3960B058186000052916442422D9600000000000",
            INIT_RAM_33 => X"9C0D46AAC79AEA56E375BA9D46A351AB526AD4B8DC6E371EA7526A000000000000000000",
            INIT_RAM_34 => X"01A2FA7D345A71D4EB6DC76C094E4511150381C0E1485659228944A2512894464E0D2874",
            INIT_RAM_35 => X"C4A2C00004600000C345A170783C1E0F078396F5EE1A94EA74E4E4395C157B31A26D2603",
            INIT_RAM_36 => X"000000000000000000000000000000000000000000000A544AAADB6DB6D874A0030D0B83",
            INIT_RAM_37 => X"A2512894462B2488945D0D568329A2B0D6ABB93ACD0EA751A8D46A351A9C6E371B8DC66A",
            INIT_RAM_38 => X"759C95634791CA16030180917D3858B2E12372476C11289D11090381C0E069365D289544",
            INIT_RAM_39 => X"8ED55A6000032F07834280188CB61B0D1800659130783C19130783EB956E0A570276DE2C",
            INIT_RAM_3A => X"D49A8D46A71B8DC69400000000000000000000000000000000000000000000086002C0DB",
            INIT_RAM_3B => X"81C0C8ED4A532D9744A25128944A231707834DAD0512B341A1D8E34E49A46EA751A8D46A",
            INIT_RAM_3C => X"EBA24E4A57038352EB329C86872390D238154280C1553459C8E52D96B6E3B12895110903",
            INIT_RAM_3D => X"0000000000052AAADB8EA6C000062113068961D1114C361B2E94D32260F0644C1E130783",
            INIT_RAM_3E => X"71B71392651A8F526A351A8D46A351AB53A9000000000000000000000000000000000000",
            INIT_RAM_3F => X"394763B1262928890381C0DB485665290ACB461118B44A25118B844532DC856B2F4ECA68"
        )
        port map (
            DO => promx9_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_11,
            RESET => reset,
            AD => promx9_inst_5_AD_i
        );

    promx9_inst_6: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"C1E0D1383E51130644C1E1458A54EA754A6575ECC68341A4DCE4ACED216860A49DC25B70",
            INIT_RAM_01 => X"0000000000000000000000000000000295606DE59180045E0F06C265A2986C465C4DA9CA",
            INIT_RAM_02 => X"42F59189CA9B67A7D36CB90AC9465A71B4A36DA8DC6E371B8CD46A000000000000000000",
            INIT_RAM_03 => X"5632D0A024E5C2E17096C8E3B13A2512888481C0CACE365D2A9485E4C2D8AC5A2316890A",
            INIT_RAM_04 => X"42A1996CB69B6D158342E1707CAA260F09842232A38A54EA74AA68B238C68F21A3CAE4F4",
            INIT_RAM_05 => X"00000000000000000000000000000000000000000000000000008BB036C0086C1E0F088B",
            INIT_RAM_06 => X"65B2E0E8562B258B44A232FA9D3E9F4FA7D3E9F4FA7D39324D291A4E27146ABEB28DC6E3",
            INIT_RAM_07 => X"71C886937754DE56B25632D8C02550B2E17096BAA3B12A251206C481C0FA63565B2E954A",
            INIT_RAM_08 => X"6DD2C0085C1911158345A29974A6D2148985616110AC22261288894352A94EA2AA7592A2",
            INIT_RAM_09 => X"49A6E351C4DE9538A3000000000000000000000000000000000000000000000000000155",
            INIT_RAM_0A => X"4540E146B55271254A65E19968C429118B8362D1390D4E9F4FA6D4E9F4FA7D3E9B51B4DA",
            INIT_RAM_0B => X"6532E94D370324949B12A71D763B24DDD538D1F69968575CB6E170B84B5B712A2510888A",
            INIT_RAM_0C => X"00000000000000010C6D8018644C1A170C8585B2D96D54561584C2E56118585A230B0AC4",
            INIT_RAM_0D => X"E9F4FA7D3E9F4FA7D3E9F4DA8DA4E55A38E4000000000000000000000000000000000000",
            INIT_RAM_0E => X"B85C1B712A2512888481C0EA6D91AA48654AA552A948565A24888542A158B446A352A7D3",
            INIT_RAM_0F => X"A230984C2A2309894AA552A954A2A92A89124E56EC89C71C884B387A32D96C6D2CB6E170",
            INIT_RAM_10 => X"00000000000000000000000000000000000089D2B124465B2C90CB65B2DA722A53098585",
            INIT_RAM_11 => X"83E1B0D86C322FA7D3E9F4FA7D36A74FA7D3E9F4FA7536D369B4DA000000000000000000",
            INIT_RAM_12 => X"7A34596CB658D2E170969CA3B13A251288C481C0E0668358D746AAA532E94CBA532996CB",
            INIT_RAM_13 => X"65D2AC6D36230A88C26130A8944612190B4AA532E94CA2AB26890A5046A4425B1D8C4B38",
            INIT_RAM_14 => X"00000000000000000000000000000000000000000000000000014A89529148C65B2D96CB",
            INIT_RAM_15 => X"4E52A954AA55298D0B65D10074445B53A7D3E9F4FA7D3E9F4FA7D3E9F4EA6D46DB6DB6A3",
            INIT_RAM_16 => X"6DB4E356312895D4F47A76996CB65B725B2D55BADB71DA2512890A81C2A06D9358D5567B",
            INIT_RAM_17 => X"6280294D16332D96CBA534D18C469B0984C26130984C24352A954AA552A94CBA23268944",
            INIT_RAM_18 => X"E9F4FA6DA6A36DB6DB000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"69A2E15D4142E8F6353DA72954AA524A954A6592188020150D17D3E9F4FA7D3E9D4DA9D3",
            INIT_RAM_1A => X"A55299707A2512894446055192BB1BA9D4F41B2B196CB65B2D57701A355B6DB85511A68C",
            INIT_RAM_1B => X"000000000000000000A5002AAD165B2D96CBA544DA7224330984C2A23098486A552A94CB",
            INIT_RAM_1C => X"45F4FA7D3E9F4FA7D3E9F4FA7D3A9F4EA6DA000000000000000000000000000000000000",
            INIT_RAM_1D => X"8E591AB1D4A111A71A71B4D3693359ECF67B3DAE9254AA552A954AA552B0D06018080544",
            INIT_RAM_1E => X"613090D4AA552A954AA532D9744A25128944A234C896412AB1E9387A1EF46CB65B2E351C",
            INIT_RAM_1F => X"0000000000000000000000000000000000000044AAACB65B2D974AA52704B196134D84C2",
            INIT_RAM_20 => X"A532E16CA8500806020180D17D3E9F4FA7D3E9F4EA7D3E9D4FA9D4000000000000000000",
            INIT_RAM_21 => X"9C2E0F7DA65B2D24CC654690ADACBC4A152BB24AEC92AD19ECF67B3D9ED75A3A552A954A",
            INIT_RAM_22 => X"242AD64C46DA3185856142E954AA552A954A65B2D9744A251289442232E88EB753AA7138",
            INIT_RAM_23 => X"00000000000000000000000000000000000000000000000000000000529B69C69B2D96CB",
            INIT_RAM_24 => X"3D9ECF67B5524A954A65D2A0A0901008040201A2EA68BA9F4FA7D46D36BA6D4E9B51A6D3",
            INIT_RAM_25 => X"A212A88AC9C09670367A4E0F67B68B2DA34AA534694CA8A30B908C590D9D8AC55CE0F67B",
            INIT_RAM_26 => X"0052936D365B2D968525AA9B7638CB0B13896132D0B4A65B2E94CB65B189544A25128944",
            INIT_RAM_27 => X"4632FACDB6DB6DB7D6000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"69CE1E8F47A3D0F67B3D9ECF67B3DAE95492A552A94850480C040201008048BE9F4FA6D3",
            INIT_RAM_29 => X"65B2A8944A25128944A251214F49C3AA70B89C3D0F67B3DB45A2D165215A74A45D2984CB",
            INIT_RAM_2A => X"00000000000000000000002AB194932D96CCEB3A84ADBA23093AC265A15974AA552996CB",
            INIT_RAM_2B => X"0100804020151117D36D34E26554EB71B8DC000000000000000000000000000000000000",
            INIT_RAM_2C => X"6D529974AA521984C265B6DE9387A4E1707B3D9ECF67B3D9ECF734D1F69974A42C141402",
            INIT_RAM_2D => X"6532D994AA552996CB65C1A0744A25128944A2511A7389C3D270F43DCE1707B3D8D5A3A3",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000295594932D96CB4C3D3614A45955B8C2",
            INIT_RAM_2F => X"5534D254A65C160A0A0100C040201008060245D4DB4DB8922D3A9D000000000000000000",
            INIT_RAM_30 => X"9C1EC6C7B3D9EF46284DC52954AA552988C261311D8F47A4E1E87B3D9ECF67B3D9ECF67B",
            INIT_RAM_31 => X"566C23360C4A74AA48664290B4A65B2D968565C1D0944A25128944A251235389C4E27138",
            INIT_RAM_32 => X"0000000000000000000000000000000000000000000000000000000000000DB4932E95D4",
            INIT_RAM_33 => X"3D9ECF67B3D9ECF67B3DAE938AC4E37197056500C0402010080402010080544A9B6BADD7",
            INIT_RAM_34 => X"A2315C7389C4E1E8B81B1EE707B3D9ECF6AA75A75AAC66332B0CC2A2511A63695CE27036",
            INIT_RAM_35 => X"00000014A68D29969B9C6A24CE06E277120A82D12954A65B2D0A8565A2D0944225128944",
            INIT_RAM_36 => X"010080402A180A888B000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"6130984DBD44AE71389C1ECF67B3D9ECF67B3D9ED74E37A2B3B40AA1D0C0402010080402",
            INIT_RAM_38 => X"65C1A064481D12894462B15C7387A4E270367A1ECE87B3D9D0F67B3A275C1146321A94C2",
            INIT_RAM_39 => X"00000000000000000000000008B42A15A8AC9C3AEC0E04EA77120A85416954A65B2C0485",
            INIT_RAM_3A => X"8982404020100804020100804020100D96CB000000000000000000000000000000000000",
            INIT_RAM_3B => X"5D581C4E2433090CC661309854A32C4DD8F47A0D4F6BA3D9ECF67B5C2E0F67BD1CE1E8AC",
            INIT_RAM_3C => X"A1A15974A04A14134382F4E064481D12074462E0C2B2B9C4E270F43D9D2E07B9C5C17534",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000C5A512137387A581C09D4EA762602",
            INIT_RAM_3E => X"3DCE1E8B83DAB270F4D1C4C1209010080402010080402010080544000000000000000000",
            INIT_RAM_3F => X"5C1D24D703A2E9D7343A3894B609230984C66122D85146236E972B7A0D948A4524D0F67B"
        )
        port map (
            DO => promx9_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_13,
            RESET => reset,
            AD => promx9_inst_6_AD_i
        );

    promx9_inst_7: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"55381C49D4EA6D96020121596CB42D0C040982C2A07038191206444560D12949C4E1E938",
            INIT_RAM_01 => X"000000000000000000000000000000000000000000000000000000000000000003515938",
            INIT_RAM_02 => X"8E2B1D756EB34E54353D9ECF7387A2E270F4560A21543010080402010080402010080403",
            INIT_RAM_03 => X"65A27064495CE360AA7A2EA4526759D24CBA75FA2C06A7144D84C24330936CB4A30984C2",
            INIT_RAM_04 => X"00000000065D5A713893275C4E04EC4D18020150F0CCBA180C068A82C2A070381D121444",
            INIT_RAM_05 => X"010080402010080402000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"61309471451E2584C2612534B1C65D1288D3954D0F67B9C3D271389C3D34615048080402",
            INIT_RAM_07 => X"4574E070381D12070365E0F95834DEC1656071EC1D49DB83AED170937A1C4A5D49A98544",
            INIT_RAM_08 => X"00000000000000000000000000025BB2713871275C4A57026D18020100E0ACAA18080692",
            INIT_RAM_09 => X"7A4E270F4D18568602010080403010080402000000000000000000000000000000000000",
            INIT_RAM_0A => X"75381C4E2351A9C6C24A309963455DC19744A225289866251289442534E55343D9ED7138",
            INIT_RAM_0B => X"01809960A42808076368A6E070381D1207064A22F2F8345A72E0E3B0476C0E0B448AE160",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000484DBD2713875371C4A54EC4D9603",
            INIT_RAM_0D => X"A251094D3520C9747B9C3D271387A3D3B415050080402010080602000000000000000000",
            INIT_RAM_0E => X"8EC76C09D6E389C760B02753BA9D4EA75313A52AD8923B84B4E494614505951855128944",
            INIT_RAM_0F => X"B86A54AE23537116020100806850180807634E292070381D120703C365F2C55C2C8936E3",
            INIT_RAM_10 => X"0000000000000000000000000000000000000000000000000000000000000DB564E270F4",
            INIT_RAM_11 => X"96C4E29D6855128944A25128944A232C2BA53A1EC6CF47A4E270ACD18541203010080402",
            INIT_RAM_12 => X"855572F96C2D66191DB04763AE070382C0E070381C0E2351A8D46AA232CE49B71DC2E170",
            INIT_RAM_13 => X"0000090A49C4E1E8F4B81A9C46A52EA627440180C04030180C149C4E5E7A90381C0E064B",
            INIT_RAM_14 => X"7A3D159DA0A8240402000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"71B09287296DC25B7096DC0E57071A528944A25128944A251089C865A5136EB953B164B2",
            INIT_RAM_16 => X"558EE4D0381A10888B8E673399C65C322555B05823ADC70381C0E0703893A9D351A8D46A",
            INIT_RAM_17 => X"00000000000000000000001B2AC7A4E2E0F4B85C0D46AD49A94ACB0180C0402010080763",
            INIT_RAM_18 => X"A25118B8442A2915134D99760365968FB415000000000000000000000000000000000000",
            INIT_RAM_19 => X"70581C49D529A8D5A93538D849BB85C2E170B85C2E170B80B1C70AA25128944A25128944",
            INIT_RAM_1A => X"AB00C040201008069CBCAD0690A81C0D88C5ACE73C1E0AAC4A2512CB3723B606E381C4E0",
            INIT_RAM_1B => X"0000000000000000000000000000000000000032EC9389C3D1D538D9DC1C6E3356A4D4E3",
            INIT_RAM_1C => X"A8D12894462D128944A251289446491307832221515136DB8E56EA000000000000000000",
            INIT_RAM_1D => X"AAB6E3B1D8EB71C5A94EA954AE2701A8D46A356A648C291CB6E170B85C2E170B84B5C6E3",
            INIT_RAM_1E => X"75DC2E0DB71B8DC6E391B4C0402010080692955E477D481C0D088BCE783399CCE44A24DB",
            INIT_RAM_1F => X"00000000000000000000000000000000000000000000000000000000369E9389C4E1D570",
            INIT_RAM_20 => X"B84B6E170B85C25AE34A250954485216894462D128944A251214852260F07832221626D5",
            INIT_RAM_21 => X"CE673399CCE44A25968EC763B60924893A6A52B88D5A9711A8D46A351A8D4A56148CE570",
            INIT_RAM_22 => X"83B7271389C4E2E0EAB85BDD6A3EA38D46E34E38D16030100806924E1ECF6A481C0E064B",
            INIT_RAM_23 => X"62B2592442260F0644000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"351A8D46A923093770B85C2E170B85C2E12D16252A30AA251088C5A231488C5A25118AC5",
            INIT_RAM_25 => X"129EE56F48540E070AACE72B3593044A2555B05823B1D8EEA648E235297526A351A8D46A",
            INIT_RAM_26 => X"000000000000000000EA3D271387A3AAE06AB83AADE68EB75BAFD469B4D3744018080492",
            INIT_RAM_27 => X"223159244221118AC5221130644221130783000000000000000000000000000000000000",
            INIT_RAM_28 => X"351AB526A351A8D46A351AB526A355BD9713395C2E170B84B6E170B84B6E094A89298A44",
            INIT_RAM_29 => X"EA34D27560100C1209B1CAD58F44DC0E070A896722555AAC4937126DC763B1DB0488D56F",
            INIT_RAM_2A => X"0000000000000000000000000000000000CB4DEC271389C2C9C66A356A752EA91C2BADD6",
            INIT_RAM_2B => X"B85C2E17096B8D295164E0F06892260C89832260F0644221110A85000000000000000000",
            INIT_RAM_2C => X"CB4763AE38E9A1B86A351AB526A356A4D5A9351A8D5A9969AA5A9BA50B25B2DB80B2E170",
            INIT_RAM_2D => X"D49AB52E371F5A15D6EA429168BA200A26094E58D58BA7542A070A69C4A25598956624E3",
            INIT_RAM_2E => X"00000000000000000000000000000000000000000000000000008A12BD270F49C3D1C6EA",
            INIT_RAM_2F => X"B8251C92DB85C2E170B85C2E170B85C2E02C96B8FAE8945214888542E1B0D8683C1D88C4",
            INIT_RAM_30 => X"6AC3225128944A24AAB05823AE371D82DF22353A8D46A351A8D46A351A8D5A9355C1D570",
            INIT_RAM_31 => X"754E27138596C2E11D351A8D5D6EB38FAD0AE4C28960385808AC094958D68B47A54E070A",
            INIT_RAM_32 => X"71A8DB693A20080402000000000000000000000000000000000000000000000000009107",
            INIT_RAM_33 => X"351A8D46A355C2E170B80B25B2396DC2E170B84B6E170B85C2E170968B25B70160B25A2C",
            INIT_RAM_34 => X"8558CF6369C68E15D38E44A25128644A256371D823B6032B8DC76F353AEE06A351A8D46A",
            INIT_RAM_35 => X"000000000003160F1AD44E154B271AC9C6A2915A0D4E385751290A8512E14C5A200A1415",
            INIT_RAM_36 => X"1636D389C51A71B69CA9A2E8803018080402000000000000000000000000000000000000",
            INIT_RAM_37 => X"B85C16570B79A8D5A9351A8D46AD49AAE170B85C2E17096DC2E170B85C2E17096DC2E170",
            INIT_RAM_38 => X"8540E070323808046804A6174F49C3D0968B4A672249C8948A25199A582C0E3B02AB60AA",
            INIT_RAM_39 => X"00000000000000000000000000000329095B12EC144AAB02A955608E9A9B86AEB42A144B",
            INIT_RAM_3A => X"B84B65A2CB85C2E170968B1475685D128803A1D100743018080402000000000000000000",
            INIT_RAM_3B => X"D43D1C6AA5538D54B2D85C2E036B83A8D46A351A8D46A356A65B70B85C2E170B85C2E170",
            INIT_RAM_3C => X"B038DC6DC35726070A81C0E070381B1005131AC4DE9389C4E149D38D44A1892D86A24512",
            INIT_RAM_3D => X"00000000000000000000000000000000000000000000062B32075B12DC24D26F4581C6E3",
            INIT_RAM_3E => X"B85C2E170B85C05970B85C2E170B85C2E02CB85C25B701628D268B8580E8944018080402",
            INIT_RAM_3F => X"3430E24D19C2CA71A88CAC964AAD43D360F49C3D164B29C2CAE16F351A8D5A9351AB5370"
        )
        port map (
            DO => promx9_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_15,
            RESET => reset,
            AD => promx9_inst_7_AD_i
        );

    promx9_inst_8: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000582CA85C31970C65C31970C6634912C964B291",
            INIT_RAM_01 => X"0000000000000000002C8000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"8CC6542914896522A1000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000004896400001428634A100000B29170C6633198CC663319",
            INIT_RAM_05 => X"000000000000000000000000000000000059000000000000000000000000000000000000",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"8CC6633198CC6633198CC64B2592CA45A319000000000000000000000000000000000000",
            INIT_RAM_08 => X"000A0000000000000000000000000000000000001349A0000050D18CC6632582C245A31A",
            INIT_RAM_09 => X"000000000000000000000000000000000000000000000000000059000000000000000000",
            INIT_RAM_0A => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"8CC65A2592CB8633198CC6633198CC6633198CA44B29850C6A3319000000000000000000",
            INIT_RAM_0C => X"0000000000000000001400000000000000000000000000000000000038C50002C3463319",
            INIT_RAM_0D => X"00000000000000000000000000000000000000000000000000000000000000000000B200",
            INIT_RAM_0E => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"8D8A000916CC663351A8C6542598CC6633198CC6633198CC66A31970A4522DA8CC663359",
            INIT_RAM_10 => X"00000000000000B200000000000000000028140000000000000000000000000000000000",
            INIT_RAM_11 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"48A45A2E18CC66B3C9000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"0016400000000000E30000143198CC66A3918CC65311A8CC6633198CC6633198CC663319",
            INIT_RAM_14 => X"00000000000000000000000000000000B2000000000000000000302C8000000000000000",
            INIT_RAM_15 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"8CC6633198CC66331948B46339A8CD6793E0000000000000000000000000000000000000",
            INIT_RAM_17 => X"2C80000000000000002C88400001400236000014233198CE47B1198CB2233198CC663319",
            INIT_RAM_18 => X"00000000000000000000000000000000000000000000000164000000000000000000B200",
            INIT_RAM_19 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"8CC66A3198CC6633198CC6633198CC6632D170C673759ACF83C1E0000000000000000000",
            INIT_RAM_1B => X"0000000000016400590000000000000000004896400000038C0059004663351E87423319",
            INIT_RAM_1C => X"000000000000000000000000000000000000000000000000000000000000000000640000",
            INIT_RAM_1D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"50C66A3D8E868233198CD4723198CC6633198CC6633198CC6632D18CF8F3519D8783C1E0",
            INIT_RAM_1F => X"000000000001680000000000000140A0005900000000000000009A2C80000008D1645059",
            INIT_RAM_20 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"F1F8EA399F0783C1D1000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"2C80000594D08450918CC6751D0D0546A319A8F6341198CC6633198CD4633198CC663351",
            INIT_RAM_23 => X"0000000000000000000000000000C8A0000000000000014000009A0000000002C001229A",
            INIT_RAM_24 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"AD46633198CC6633DAED76A33D1F0783C199000000000000000000000000000000000000",
            INIT_RAM_26 => X"0000000002C001B6914C000011A4C06CB2D18CE83A1D8A8C663359EC74233198CC663319",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000002C800000000000005900000B200",
            INIT_RAM_28 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"E868233198CC663359CD46633198CC6735E3F1D6793E0F0783C151000000000000000000",
            INIT_RAM_2A => X"00000500000001340000000000070284B4984C001B6E04890CB519C8EA7B1A88CC6723D8",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000002C8000000",
            INIT_RAM_2C => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"C8EA7B1918CE47B1D8E868233198CC66B3BB8CC6633198CD6BC7E3F1D47C1E0F07833319",
            INIT_RAM_2E => X"0000000002C8000000000A050280000134000000000006845530E02C245B2E010890B322",
            INIT_RAM_2F => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"F1D67C1E0F0782A319000000000000000000000000000000000000000000000000000000",
            INIT_RAM_31 => X"0036DC09821891A3A9E8743B119A8F4343D0EC54633198CC67C79A8CC6633198CF8FB5E3",
            INIT_RAM_32 => X"0000000000000000000000000002C8000000000C000590016450002C00000989126930E0",
            INIT_RAM_33 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"8CC663319CD78FC7E3E5747C1E0F0726A351000000000000000000000000000000000000",
            INIT_RAM_35 => X"2C00000E0DA161A0D06D261C0590E06AA3A8E87634119EC763B5D0EC46633198CF8FC719",
            INIT_RAM_36 => X"000000000000000000000000000000000000000000019108000000140000091002680098",
            INIT_RAM_37 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"EC4663319CD78F95198CC663351F1F8FC7E3E5783C1E0F066633C9000000000000000000",
            INIT_RAM_39 => X"2C800005900268B0980000131228D440B298A1B81C0230E26B25D0EC762A3A0E876395C9",
            INIT_RAM_3A => X"000000000000000000000000000000000000000000000000000000000000059140000000",
            INIT_RAM_3B => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"E87635199E874393DAD44663351F1F8EB519A8C66339AED78FC7E3D4F83C1E0E8D4761D1",
            INIT_RAM_3D => X"0000000590000000300000134000036A205800161C19E48A60B5224C440B2434A38F53D8",
            INIT_RAM_3E => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"D5783C1E0E8E67C1D2000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => promx9_inst_8_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_1,
            RESET => reset,
            AD => promx9_inst_8_AD_i
        );

    promx9_inst_9: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"70260241C4DEABB1D8EC74351DAE876393E3A8C6633E3F1F8E33198CC6633E3F1F8FC7E3",
            INIT_RAM_01 => X"00000000000000000000000005A0000000500000134002CC65C0000038232A48CA84435A",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"8CC6735E3F1F8FC7E3E4F83C1E0F0783A3E3000000000000000000000000000000000000",
            INIT_RAM_04 => X"4C382A65A7004936E07016848658D6A3B1D8E8763A1E4D4683B1E4A8C66B3E3F1F2A3319",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000590000050500000122586D381C000",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"70C67C7E3ED66A33198CCC3B5E3F1F8FB5E3E9783C1E0F0783C7E3000000000000000000",
            INIT_RAM_08 => X"0000244586D3813058702622A9A54869B6E04C06D7ADDC8D67A1D8E8743A1ECEC72B93EC",
            INIT_RAM_09 => X"00000000000000000000000000000000000000000000000000000000000005A000005000",
            INIT_RAM_0A => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"EC763A1EDEC78F93ED9856BB5E3F1E8633198CC8BC7E3F1F8FC7E3D4F83C1E0F074BC7E3",
            INIT_RAM_0C => X"00000005900000B2000016244008CB81C0E07048835222C98DB2E02D06D391BACE87B1D0",
            INIT_RAM_0D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"E9783C1E0E4F8FC7E3000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"09375889A6D763B1D8EC763B1EDE4EEF43ED70F8FB5E3F1C6633598CF2BC7E3ED78FC7E3",
            INIT_RAM_10 => X"00000000000000000000000005A00000A0002C3824458AD381C0E07037086D92D26CB2A1",
            INIT_RAM_11 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"8CF8FC7E3F1F8FC7E3E4F83C1D1F1F8FC7E3000000000000000000000000000000000000",
            INIT_RAM_13 => X"4C37138980D310B21211B753ADBACF63A1D8E876395EDE4FB3A7EDA8F8FC7E3ED466339A",
            INIT_RAM_14 => X"00000000000000000000000000000000000000000005900160B0004C3824498AD381C110",
            INIT_RAM_15 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"ACF8FB5E3ED387359AAD78FC7E3F1F8FB5E3F0783A3E3F1F8FC7D1000000000000000000",
            INIT_RAM_17 => X"7038244D0AD381C0E06DA6D36A14E08C241B6EB704654E8763B1D8EC727B5EDD0FB735EC",
            INIT_RAM_18 => X"00000000000000000000000000000000000000000000000000000000000005A00160A058",
            INIT_RAM_19 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"F26A3C7ECE9FB3C99CED78FB5E3CD547C791F1F6BC7E3F1F8FC7DAF0783A5E3F1F8FC7D1",
            INIT_RAM_1B => X"00000001914260609870382B519882615298AA06938594D84824236EA7418DBD0683B1D0",
            INIT_RAM_1C => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"F074BC7E3F1F8FA5E3000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"6E0301959ACE83B1CAED743D9DDF2793C9E3F1F8FC7E4CD78F779AF1F8FC7E3F1F8FC7C9",
            INIT_RAM_1F => X"0000000000000000000000130282CA60A11070382B55A70285A098AA98C34196204836DD",
            INIT_RAM_20 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"F1F8FC7E3F1F8FC7D2E4F6FC7E3F1F8FC7E3000000000000000000000000000000000000",
            INIT_RAM_22 => X"8AB10345A4A84848DD4E87039A091763A1ECE5727DBECF67B3D9E4F1F8FC7E3ED78FC9DA",
            INIT_RAM_23 => X"00000000000000000000000000000000000000001C0002D380B0E070382A75A4C169C05A",
            INIT_RAM_24 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"F1F8FC9E4F1F8FC7E3F1F8FC7E3F1F8FC7C9E9F6FC7E3F1F8FC7E3000000000000000000",
            INIT_RAM_26 => X"70382455328169C09B4DA6C249B118713ADC0E030B6DBACF6395EDE4F6BC9ECCDFB3D9E3",
            INIT_RAM_27 => X"00000000000000000000000000000000000000000000000000000000161C0002D3813110",
            INIT_RAM_28 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"D4793D9EDCDFB3DBDAF1F6BDBE3ED7B7C7E3F278FC7E3F1F6BA7DBE9F8FC7E3F1F8FC7E3",
            INIT_RAM_2A => X"0026220002D38130E070382B5221096522DC4DA6C36AC06031B8DD0603136B3E8683D9ED",
            INIT_RAM_2B => X"000000000000000000000000000000000000000000000000000000000000058000013000",
            INIT_RAM_2C => X"E9F8FC7E3F1F8FC7DC000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0603136DBEC72BD9EDD07B7C9E3CD7B3D9DAF1F93D9E3F1FB3B5E4F1F8FC7E3ED78F55D3",
            INIT_RAM_2E => X"00000B0DA00001520000261C0582CB81A0E070382332209164B2DC2D2703494061722A1C",
            INIT_RAM_2F => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_30 => X"F1F8FC7DAF1F8FA7E3EDF4FC7E3F1F8FC7E5000000000000000000000000000000000000",
            INIT_RAM_31 => X"2D98C349506311580C0E0303959E87B3D99CCD7B3DB91F6FB3C9E3F1FB3D9DAF2793B5EC",
            INIT_RAM_32 => X"00000000000000000000000B35A00001C05800381C0982CB8190E070382331309244B55D",
            INIT_RAM_33 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_34 => X"F27B3C9E3F678FC9ECED78FC7E3F1F8FB5D3F1F53C7E3F1F73CBE5000000000000000000",
            INIT_RAM_35 => X"8844244DB0D164259E4D869581C0E3753A1C06030A9D8E57B337E4F67B3C7A0F6F93C7E3",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000123DA2C002205800441C0E000365A0E0",
            INIT_RAM_37 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_38 => X"F67B395CAF67B7C7E3F67B377ECEEF6BC9E4ED78FC7E3F1F8FC7D3EA753C7E3F1F97CBE5",
            INIT_RAM_39 => X"00381C0E000269A0D070382B4DB0D164355D4D849361C32C54380C0603137D8DDFB735EC",
            INIT_RAM_3A => X"0000000000000000000000000000000000000000000000000000000C8A135E39800240E0",
            INIT_RAM_3B => X"F6753C7E3F2F97CBE5000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3C => X"0603245A1F679393ECF67B351DDF678FC7EDF6793C9ECF278FD9E4F1F8FC7DAF1F8FA7DB",
            INIT_RAM_3D => X"0C884B7E3E4A6261504C38220E04C285C0D07038244DC0D048C6DC4D869360C4E270180C",
            INIT_RAM_3E => X"00000000000000000000000000000000000000000000000000000000000000000000B600",
            INIT_RAM_3F => X"ED78FC7EDF1F4FA7D4F278FB9E5F2F97CBE5000000000000000000000000000000000000"
        )
        port map (
            DO => promx9_inst_9_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_3,
            RESET => reset,
            AD => promx9_inst_9_AD_i
        );

    promx9_inst_10: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"4D869380C8A994381C06072B35BF672B37ECF276B93ECF6F6BD9ECF6793D9E4F1FB3D9DA",
            INIT_RAM_01 => X"10800000000164325C0906C25E3E56A131A97044220E070165309870381535D0D04936DC",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"F67B3D9E4F27B3D9E3F1FB3DBE3F1EABC9ECEDF73CBE5F2F97CBE5000000000000000000",
            INIT_RAM_04 => X"70441315D21848C6A44D8693A24AF090180C06152B3EDF6CC3D9ECF6F43B5E4DDF93D9EC",
            INIT_RAM_05 => X"0000000000000000280C884425A0016C361B2D8B027D3F1F62B3D08854240E088261A2D0",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"ED6A3C9ECF27B3D9ECF67B3D9E4F67B3C7E3EEFB7C7E3E9F53D9D4F2F97CBE5F2F97CBE5",
            INIT_RAM_08 => X"E838350E07038142D070380B2DC3190CC6DB4D86D2A956E030180C0626E57DDCD647D9EC",
            INIT_RAM_09 => X"00000000000000000000000000000000500010970005C0C88428140A06DBB1BF1F2BB1D0",
            INIT_RAM_0A => X"F2F97CBE5F2F97CBDE000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"0616E795CD0F2BD9EDE4F63DBECF67B3D9ECF67B3C9E4F279377ECF678FC7D3EEFB33BE5",
            INIT_RAM_0C => X"16455B934F1F8FB1D0EC743A0E07044134E068380B2DC4D97136DC4D90CB8DC4E870180C",
            INIT_RAM_0D => X"00000000000000000000000000000000000000000A0000006432122D86C5812160482814",
            INIT_RAM_0E => X"DDF4FC7ECF2753AB9EF2F97CAD5EF7964C5A000000000000000000000000000000000000",
            INIT_RAM_0F => X"4DAB0393E21830180C06172B9ECE878FC9E3E872BC9ECF67B3D9ECF67B3C9ECF27B3C9EC",
            INIT_RAM_10 => X"09394362C0A05028140A4D3399CF1F6BC7D0E8743A1598CB81A0D94844122A49A274B934",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000000000000000016400D110800B25B",
            INIT_RAM_12 => X"F2793D9ECF67B3D9E4ED793D99CCDF5AAB55F2E794B9EF2B70279E000000000000000000",
            INIT_RAM_13 => X"70380B49C8E9716C9B52370493406090380C1236F35DAD4793DBC9E878F37ECF6793D9EC",
            INIT_RAM_14 => X"5080142284D16424124E9714A1C0A05028140A173DBA5F676BC7C9E8763A192A8B81C09A",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000980000000000000000000000000A1",
            INIT_RAM_16 => X"D466BDBECF67B3D9ECF67B3D9ECF67B3C9E3F67B3C792EB455ABE5CF2962BDE4E0728DE5",
            INIT_RAM_17 => X"D0763A154CDD66A29A6838166A58A9716D1D4E270471D1209018246D743A7C9EC7B7C7D0",
            INIT_RAM_18 => X"00000000000064500070B8530918D048245A2E2D16C9D0E05028140A29269E4F67B3C7E3",
            INIT_RAM_19 => X"52B573C5C0A273CBE50000000000000000000000000000000000002C0000119000000000",
            INIT_RAM_1A => X"E8763C7D0E57B793D8E4F2BD9ECF67B3D9ECF67B3D9ECF67B3C9ECEEF6B33D6AAADAAB9E",
            INIT_RAM_1B => X"0E33669DDAD7B7C9E3F1F435359AAD6BB910A9C65B4B6932916CC67297098CD2609048E3",
            INIT_RAM_1C => X"0026001506800000000000000000016232E148C65A31964168245C0DB596CB65B0702814",
            INIT_RAM_1D => X"E56A7AB5563357BCD55B519381409F5BCBE5000000000000000000000000000000000058",
            INIT_RAM_1E => X"630719A2C1613059A0E874333D0E578FA1D0D066FD9E4F2777D9ECF6673D9ECF2793D9EC",
            INIT_RAM_1F => X"4EAD96CD58AB18CA1C4E16A69E4F646BD9E3F1F2753AA8E773C79AA968966C65B2756CB6",
            INIT_RAM_20 => X"000000000000000091004640150A88000000000000000140A0B1198CC65B3198CB68365A",
            INIT_RAM_21 => X"F666BC9ECF67B3D9CAD47733CD56351AAAB66AC543814AAF97CBE5000000000000000000",
            INIT_RAM_22 => X"AD78DB2C66B2D98CC6632946A2C0A0B0B5D0E874393D0F66A3B1D8EC7B7D9ECF678F77DD",
            INIT_RAM_23 => X"8CD6D90E18CC64245C4EB196CB68AE7298DC4E66D67A595C8BD9ECED78F234389D57C7DC",
            INIT_RAM_24 => X"000000000000000000000000000000000059884823351E4A60000000000005900345A2C8",
            INIT_RAM_25 => X"E4FB7C9EDDDE47DBECD0FB3D9ECF67B337D0E97962AB66AE796CB69304C285CEF797CBE5",
            INIT_RAM_26 => X"F278F39136AB57C7E3F1F73B6D55B4F96D466AD186A140A0513791E8763A1D0ED763B1D8",
            INIT_RAM_27 => X"0036400006880235198CC8BDAE14C365B51D4EAD96CB66AD57B9DCCE773B8DA95B6933ED",
            INIT_RAM_28 => X"2E050294CF2F97BD55000000000000000000000000000000000098A8D47C1A1E95440000",
            INIT_RAM_29 => X"EC763A1C9D0763A1D8ED7B3D9DAD478FC9E3CD7B3D9DDF2793A1D0EAF794AB6A34556CD5",
            INIT_RAM_2A => X"CE78FC722ADA613122F6F8F37156AD33C7E3F1F8F39156ACD98D9E8AF9CCA5C6E170291A",
            INIT_RAM_2B => X"68727A3E0E9781300000341300048A8523198CC6735E691261409A933556CD6CF51AABDC",
            INIT_RAM_2C => X"F2B556CB68AAD96CD50A050B9DEEF5562B550000000000000000000000000000000000D9",
            INIT_RAM_2D => X"A379D8D15AB2B028DBCD68393A8E4F43B1D0F1FB343D0D47B7C9A8F2777D9DDCAEA3A192",
            INIT_RAM_2E => X"4D49B3D46CF79FCFDECF77BB95A4C3693090ADF7738D58AE8BA5E3F1F722B3E6ACDB3D46",
            INIT_RAM_2F => X"000000000000000058E4D4393D2E974BA25800263325948465C3198CC66339CF636530E1",
            INIT_RAM_30 => X"F27B3C934E9F43A1D5F2AD96CB6632D98C350A051ABD56AB59CA1C000000000000000000",
            INIT_RAM_31 => X"F1E76694F8F47B7DE7F3F9F3D9EF32919AE3CDF2795CAE4E87B1D0F6E87B1D0F1F9341C9",
            INIT_RAM_32 => X"8CC663319F6FB1C2A04C4733DE7F3F9FCFE7EF79FCB224C26140D92C56DCAD68E683A5D2",
            INIT_RAM_33 => X"000000000000000000000000000000000000A854741E3E8F8FA39900163535968B463319",
            INIT_RAM_34 => X"D0F63B1C9F6683A1BBF27934AE5D474353E58AAD96CB6632D96C1C0A0524CA5631702814",
            INIT_RAM_35 => X"AEB718CB6D1783A5DCF1F8F6D4E9BCDF3D9EF3F9F3D9EF3375BB1BCE66B779BD0F27B5D0",
            INIT_RAM_36 => X"CC8033359D846633198CC66B4E1ADF9348904C242DDE7F3F9FCFE7F3F9FCF9C8CA653098",
            INIT_RAM_37 => X"0E2956CB60E05028B400000000000000000000000000000000000068783A3D2F1F8FB7E0",
            INIT_RAM_38 => X"D2EEF39ECCDE6B95D0EC763A1BBD474393ECF6F75AB13E8763B9E55B2D96CB65B2D8CA14",
            INIT_RAM_39 => X"F3F9FCFE7DF26930A06D6794B4CD1747A5D4F1F7337958F2919B56DF79FCF9ED2E9438AC",
            INIT_RAM_3A => X"2C727A5D2F1F8FC7D2F06676130ACCC233198CC66459C70FB3D92B4C28239E7F3F9FCFE7",
            INIT_RAM_3B => X"5B2D96CB6633186A1C4EAD96C1C0A0506B260000000000000000002C8000000000000000",
            INIT_RAM_3C => X"CF79FCF9EF34D85823D2FB7D9ECCE7B351DAD468741D0E8743C9ECEEB958D92EC743AB55",
            INIT_RAM_3D => X"4C281A3E7F3EFA389A2CACEABE7F3F9D429868F9D8D9AD0F47A5D4EA753C9DD4DE7AAAC4",
            INIT_RAM_3E => X"09064000000000B0D90068743D2F1F8FC7DBF06C393A98CD4633198CC66B75ADDD6FD9ED",
            INIT_RAM_3F => X"8AADA39D0EC64BCAD55B2D96CB65B31838A55B3186A140A071ACB6000000000000000000"
        )
        port map (
            DO => promx9_inst_10_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_5,
            RESET => reset,
            AD => promx9_inst_10_AD_i
        );

    promx9_inst_11: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F6F53BBED8F533CB9BACC8ABB5C6E17046946DFB3D9E4F656B779AED727B1D0E872BD9DD",
            INIT_RAM_01 => X"8CC66339CCE7B3D9ECADA80B1BE5980000122D8483259F3F9F3C686DF9E8DD2E4D47C7D3",
            INIT_RAM_02 => X"0000000000000000000C88400000000001A188383A5D2E978FC79AE9E82B3998CC663319",
            INIT_RAM_03 => X"CD743B1D8E87B354DC5B2DAB5D0E8772AAB6632D96CB65B2D94AB65B19428140E2D96CB6",
            INIT_RAM_04 => X"AAF9E8DA08866E9913CE7B7DBE66E677CBD4D0C654200000A12A668F57279E4F67B735D3",
            INIT_RAM_05 => X"8CF4F5359A8C6633198CC66455AEEF93C9ECF6A4130910006CB8140A0B028122C79FCEDA",
            INIT_RAM_06 => X"5287028355B2D96CB6000000000000000000090480000000A0B0D0E8C83C7D2F1F8FC7DC",
            INIT_RAM_07 => X"2A1957BA5F27B3D9E3D4763A1D8E4D663AC65B45751D0D4F59AAB4632D96CB65B3196CB6",
            INIT_RAM_08 => X"0C864362C0944FCF4CCF79F43C954ACC245A2D673DBE6F379B3B9AE8646329800558CA66",
            INIT_RAM_09 => X"E9683A5E3D178FC7E3ACC66B319A8C6633198CC66B59BCDFB3D9ECF246CB0282D86C2412",
            INIT_RAM_0A => X"6AAD96CB65B2D96CB61A850CAC65B2D98D460000000000000000000904C000000001C658",
            INIT_RAM_0B => X"E8741C2988DD3A6EE633198AA54D2CF3DB9BF1E87A1D0AD4554AC66AD6723D0EDD562ADC",
            INIT_RAM_0C => X"F67B400000C848241209048241316003CF9EF3F5B42980904836A48DFB7CDE6F37B7CDD5",
            INIT_RAM_0D => X"0D86C00000000138D9A874BA5E3E978FC7E3E9C6633518CC6632E18CC66335BF67B3D9EC",
            INIT_RAM_0E => X"A9D66A9A8EB396B315632D96CB65B2D96CA50E0D56CB65B2D9ABD6000000000000000000",
            INIT_RAM_0F => X"D27B3CDE6F379BCDD6D4B2000DADB4DDCC6E33198CC0C2E36FDBE4CE66AB51C6AAD96CB6",
            INIT_RAM_10 => X"8CB86B4E1CE7B3D9ECF67B1B4280008424120908424120A04B3DE7F3E6A2000090B098DC",
            INIT_RAM_11 => X"00000000000000000016050001900160B92BA874BA39BEE78FC7E3F1D6AA3198CC66B559",
            INIT_RAM_12 => X"2D8516CB6632D96CE5AD457259B8AD6AB4B65B2D96CB65B2D98C350E2D96CB65B2DB3C9C",
            INIT_RAM_13 => X"F3D4400210D86C3995F27B7CDE6F379BCCDAE4C81B5EDA7CDE6F4F93258CC660E49A7934",
            INIT_RAM_14 => X"F1F6DC3198CC65C39B70D6AB55B8CFB3D9ECF67B34A001406424210004858140A04A39E7",
            INIT_RAM_15 => X"5B2D96CC65B499381C0000000000000000210A06CB20014000B896CCF4BA5A2CDF8F37E3",
            INIT_RAM_16 => X"4A198CC351E95269346E050CA9D5B2D98D1372C7353B4AD6A5CAB65B2D96CB65B3194A1C",
            INIT_RAM_17 => X"0905028140A04A27E78A8A000120D850B934F6793CDB6F36DBCC59E84C1B5A59BD3E6EBB",
            INIT_RAM_18 => X"6EE83C7DC68772B59BF1F8EB5198CC66335ACE466B79BCE56FD9E4F2793DADA0C8A00000",
            INIT_RAM_19 => X"5B2D96CB65B318B8B6633196CB66B270380C0000000000000000120A04C24190C864CC66",
            INIT_RAM_1A => X"4C546B7A4A74DE6F4F8DA74CC6633070985C0E050CAA552AD96CC66B6479359D4D4D6CCE",
            INIT_RAM_1B => X"F667349A50C86450DA2D850281B0904A391C18250241B0A0B34BECF279BCD1EDB39A4C94",
            INIT_RAM_1C => X"0A04836212C8852C663346F33E38D467B8D9E9F8FB9308CC66B4E1CE66E359CCDFB3D9EC",
            INIT_RAM_1D => X"AD762B3AA8D3193B575B2D96CB65B2D94AB6633198CC662070183D00000000000000001B",
            INIT_RAM_1E => X"CAEAA78E632C98AA664A26337A5A753E6F4FDB67A6C6533198582C0E0506A5C5B2D96CC6",
            INIT_RAM_1F => X"8CEEFC99BF66EFD9ECF67B542BB9A06434285606C24120904800191E86836140DE97D9D4",
            INIT_RAM_20 => X"00000000000000005C0A048285A0C88D2C653325A37E3ED9A2B59B6876FC79B8CC6633ED",
            INIT_RAM_21 => X"5B194CAA55B2D98D13CCC4EAB138AA963CCE5B2D96CB65B2D9AAD5632D96C4C0603048AC",
            INIT_RAM_22 => X"2D06858146E657A7E3EA6A64C9633258CC663316AB756A74DE9D379E48BAB5E5F170281C",
            INIT_RAM_23 => X"6D287A7DC8CC66335BF6E73D9EDF27B3D99CEEF9256590D068745A00064241210864C65C",
            INIT_RAM_24 => X"63318FC1C0E2522AC600000000000000322C0A0486A5B091712C4C2A90DB71BCDC693192",
            INIT_RAM_25 => X"A7CAEA73E5F1B8982C0E3196CB65B2D96D1C8AB95B9155B4DA9EB6633198CB66AC564CB6",
            INIT_RAM_26 => X"2A16850212C96834210908C58146EC4FC7DCF1EA2B69633150CC553316A57ED9BCDE9F37",
            INIT_RAM_27 => X"3B131B4DA95F4D2090AD3852192E9C6632E1F27B3C9ECF67B3C9E44D4D268212A030380C",
            INIT_RAM_28 => X"5B2D9AB26932D96CB65B274485C6EA756CB600000000000000425C1A848B81B0906CCA4C",
            INIT_RAM_29 => X"4B0A3DB4EA7CDE9E5A9353E379C6E998984C0A1956CC65B3568D15633962ACE9B53E3CB6",
            INIT_RAM_2A => X"F6964341C06030380C0E0303854118E824120908C58144E66FC7D2F1F43A0DB33048CC5C",
            INIT_RAM_2B => X"3284CCA1416048984C161D937195DB6AB4984C369C2908D751919B8CD6FD9ECF6673DBED",
            INIT_RAM_2C => X"52CDA6D569BCDDACB663456BCC65B3196CB663131BA9C4EB196CC6000A00000000002414",
            INIT_RAM_2D => X"EDF43A1514A86CA8232E46FBBA5A74DDCCDD31D3E6DB4CF374CA140A0D54AD5A34556CC6",
            INIT_RAM_2E => X"ADFB7C9ECF6570B09A2C8E8B654118E846231186C361B0D86C241B0916CB65B8E78FC7D2",
            INIT_RAM_2F => X"0016400000016836351A8D4CA140E06C287E16130595ACD322331A4C26130A14C24234D1",
            INIT_RAM_30 => X"2E3962AE56AB55AB3EABC7A3D4FA7CDA2B268ACD99CC66B359AB268AA50989D632D96CB6",
            INIT_RAM_31 => X"09366B359CDF73B792D4F43B0D92D06CB812096572BDDD2EDA9E63623999DDEEF3752C76",
            INIT_RAM_32 => X"8CA6140984C28130C84C242575CD24F1CC5B0E070A8301086836120906C361B0D8483612",
            INIT_RAM_33 => X"121316CB65B2D96CB6001683230000B036650E194CA351A850382C1A93028DAF1EED9099",
            INIT_RAM_34 => X"2DD3E9D55F2B7588CD72A722B269F67AAD57ABD5EAD5EAF4996CB69B4D94AE59F49A4C9C",
            INIT_RAM_35 => X"0904824120906C241209168D3A0D4F8FC7A9D4F43B0D90D84836122649B2B95D26966EB3",
            INIT_RAM_36 => X"1A850289BCCF6B76C84C26140A15028130A0501A540692187038542A084605818068741B",
            INIT_RAM_37 => X"AF49A7D9E6AAD898243F3196CC65B2D96C246D54CC69A4D8506A651AA746AA5328702835",
            INIT_RAM_38 => X"262DB2AE5F6F774BB60D47A6F9EF2E397CCDAAC763B5DCF55B3D56AB55AAD578EAD9AB36",
            INIT_RAM_39 => X"18160B0582C86824120D848361B0D848361B0D969B519C8F6FB7D0D4F63A119090484623",
            INIT_RAM_3A => X"52B1838C632994286532850285BACF8FB5E370A6140984C26130A15096C74430E0307421",
            INIT_RAM_3B => X"AB55AAD5E8ECFABD5E6755A9ECE6B13098B65B2D96CB65B358984C50C4C46590C8B1381C",
            INIT_RAM_3C => X"E874341191D08C461C262D9CAD68AE71B9ED9E18F6C94CF7962ADC6D465B3198CB69B756",
            INIT_RAM_3D => X"4C280B6540603086582C0A130911808424120D86C24120906C2412090693519A8F4B93A9",
            INIT_RAM_3E => X"0D064A81A10850B89C5B194CAB65B294286532850281B8CF6BC7BBCD3693098502614298",
            INIT_RAM_3F => X"8D54EA753ADE974B56AB55AACCEABD5DBD36934DE6CB6329F98CB6632D96CB65B130495E"
        )
        port map (
            DO => promx9_inst_11_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_7,
            RESET => reset,
            AD => promx9_inst_11_AD_i
        );

    promx9_inst_12: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"1D369B3198CE4755D0EC742B29A091501823262D96CD55B47549A5CE57279E6AEF97CB9D",
            INIT_RAM_01 => X"8CB2130A05028130A050A60D021109A442589174F545810848B43A0906C241B0D8483612",
            INIT_RAM_02 => X"5B3598CB6260912C9C1086446120C85028B452B194A655B31838A532850282C6D56BB551",
            INIT_RAM_03 => X"F6B8FBBECAE67BCBD58D46633198CCD1BB4EA74DE9F379BC7A9F379BD3D4A9D5B2D98CB6",
            INIT_RAM_04 => X"09048241B09048365A6CC6633518CD4751D0A8D6740A10908C181C0E2D96CB663356BADC",
            INIT_RAM_05 => X"328D4285C6D46735E3F1F8F34E14C26140984C28130682C14233D3F1F70B2914D469421A",
            INIT_RAM_06 => X"9BAD96CC64EB39ACB6673596C7E0E03038650D884241C1086C289CA62D98C9D5B2D8CAB6",
            INIT_RAM_07 => X"329316CB6632DA4DECF637269ECD24D3CBE5EAB4633198CB6668BD934DE6F379BCDE6F37",
            INIT_RAM_08 => X"EDC67355AACB40421B0906C34120906CB4D98CC6633198CC663391D0285349A0908C863A",
            INIT_RAM_09 => X"A6355AA655B2D98C6563194B65B4D46735DAF1F8FC7BBCD46530984828520304C56BB9E3",
            INIT_RAM_0A => X"A753E6F379BCDE6F4F9F2D94ACEAB2F96CCE9F2D8981C06091CC652A084341C090682814",
            INIT_RAM_0B => X"64364D25A4D9A4746856131ACB65B319CB34F6774B7ECF6573ABE5F2E6E33198CD6F4BB6",
            INIT_RAM_0C => X"ADA40A159E978FC7E3F1F6F43994C0C03612090C024124D049B3198CC66331A645723319",
            INIT_RAM_0D => X"0E04832232A064365B89D556CD55B2D96CB663194B65B6D46735E3F1F8FC722ADEEF779A",
            INIT_RAM_0E => X"F2F5769538CC65431B5DD3A6F4F9BCDE6EE64ECFA9F269B2DA6D575B130181C2A4DCB81C",
            INIT_RAM_0F => X"8CC663322A747A9F4FDB26130984C28540DA2D2D8FCB65B2DA3ADCCE7932BDDEEFB559E5",
            INIT_RAM_10 => X"F1F8F375B09169345A10A6B33A0EDF8FA5E3F1F839298180E8365A18164B4A16CA6A3319",
            INIT_RAM_11 => X"26090B8E6ABA50B91E1207034120E068285A2D7722AB6632D96CB65B318389A6D385C39A",
            INIT_RAM_12 => X"ADFB2B99CF6792B9E5F2D4F37B4DA5533943D2D5AAD56AB53A9D57ABD3E6F3672CDAAE9D",
            INIT_RAM_13 => X"2C9A533196CC6633198CC65C32BA7D3E6F4F4CA6142A04C264B29072AD8CAB65B2D9AB9C",
            INIT_RAM_14 => X"5B354CADA71C663319ED78DB7BB2D0E824122D567A3D2E9687C7D2F072530300D8686058",
            INIT_RAM_15 => X"CF57A7D6EAF55A6D1D6EC7AAD3466C56AD5E0910C741A11870345A2D68B399C8AB556CD5",
            INIT_RAM_16 => X"4DB196CB65B2D96D1DCE7B7DB9DEA777BBD6F2E6E3319A1C4EA79ECF67B3D9ECF63B3D9E",
            INIT_RAM_17 => X"E8B40B05A108C0B0A12824233198CC6633198CD46574F9BCDE6EBB8CA6130A04C345B89A",
            INIT_RAM_18 => X"2D467B9DC8AE716D155B295CA9B4D46632BB70C8A78B36D84836126D467A3E0E978F43E0",
            INIT_RAM_19 => X"CAD5ABD5ECF67ABD9EAF576BD5EAF57948DDAB55AACDD8F55AAD364D048363A0D070242C",
            INIT_RAM_1A => X"EA261A0984CA6D38B65A3196CC65B2D96CB68DE6FC95DCEF53BBD5A954EB7438CD6A34DA",
            INIT_RAM_1B => X"4D667A3D2F1F4BA5E09016042301824232C88CC6633198CC6633198CB869F379BD3E3C98",
            INIT_RAM_1C => X"CE268361B1D08C481A2D383B9E3F1F722B9C8AB55B4A46D38632DA2A26CB60C2A1503612",
            INIT_RAM_1D => X"A1B69A31AA9D4EA75B6455A9F57AB55AAD36AB55AADB68F376AF578F271BB4FAB55E4CC4",
            INIT_RAM_1E => X"8CCD26F379BD3DA3D4CDF4F389871A95CAB65B2D96CB65B2D96CB68EF8FD9DD8AF53A9D4",
            INIT_RAM_1F => X"21870180C1186C245ACCE83A3E3EDF4BC15128160B02170C6633198CC6634E18CC663319",
            INIT_RAM_20 => X"6F53E6F4F9BCDC4854DF67136120D86C861A11B82A5E3F1F8F399C8AB5634DA8CB86449A",
            INIT_RAM_21 => X"6ACC349E4CAF77A9D4EA46D36544DA69B553CACD2AD57A74DEAF4FAB55AAD56AB55AACDD",
            INIT_RAM_22 => X"6D268B3198CC6633198CD3A6F37A7D6FA722CD78DB31359AD96CB65B2D96CB65B3196CA5",
            INIT_RAM_23 => X"CE671CB198CC66325421830180C0E06C2519ACE87B7E3E974792982C140249A70B6A329A",
            INIT_RAM_24 => X"A7CDE9F4EABD3EAD56AB55ABD5EAB270B8244C553A89A71848341B0D26AA3E3F1F8FC7DC",
            INIT_RAM_25 => X"5B2D98CB65B2D96C655B56AB3EDF666F39D4A1C69BADD2E09128DA9A38F6D56AB57AAD56",
            INIT_RAM_26 => X"1808D369A2E268B4120904935198CC6A33198CD3E6F4ED2E6FB891EE797ADD5EAB556CB6",
            INIT_RAM_27 => X"0D08DC1DCF1F8FB9A2EE773391A8CC66325B0603018231186DB49ACCF4BC79AE9745B258",
            INIT_RAM_28 => X"6ECF24D4FABD3E9D56AF57AAD56ABD5E9F26A753E9D264A195BB1E14161B5B4CDD0DC612",
            INIT_RAM_29 => X"EE797CBDEF2C722AB65B2D9AAB65B2D96CB60E397435BF6753C7D4A1B6934244EB75BB57",
            INIT_RAM_2A => X"E8F8FB7D2F0684B02816050582C0A06C46120904A3319AA56A459B9A53AAD4F8D74C0152",
            INIT_RAM_2B => X"000A0B0506D7733743118693519CD66BC79BF1F6F359B8CC6633192A030381C0606CB559",
            INIT_RAM_2C => X"CD54D765406070B8C48F55A9F4F9BD3E6F37A7D3EAF56AB47A6D36AB55DBC4C4A499CC24",
            INIT_RAM_2D => X"DB55B492B4D000019BDA797CB9EA6639B34C6AC56A515632D96CB632A76355ADDF53A9DA",
            INIT_RAM_2E => X"2D830180C0D84935E0CD74BA3E0E8A60505C0A05028140E06C24120955339D5AD54FAAD9",
            INIT_RAM_2F => X"8F312AD56AB375386500000000028162A7DCCDA703691CDC67B79AA974B355AAD54632D9",
            INIT_RAM_30 => X"52871C79BAD6EFC7D49146588AC12070381C12251BB1EAB47A3D579BCDE4CE64B39A9F57",
            INIT_RAM_31 => X"09473CBE5EB79737D4ADE974A980000000A9A9F5BAD6ECF370B5508AD4AA5518AAD96CB6",
            INIT_RAM_32 => X"ACE6EB519AD465B29B0E150181C0904AB3E0E4F83A3E0A8960B6120A050281409048251C",
            INIT_RAM_33 => X"6F258CAE69BCDE6F269BCDE6E95120712A6E000000000181405050A9F73389C54C81C152",
            INIT_RAM_34 => X"D0D4B35E0D13194AB65B0D5B922AD76BC7D3CE18CB6946E970380C1A8D47A5C4EC7A3D1E",
            INIT_RAM_35 => X"0A05036120904938DCAAF97CBE5F2F9739D4F6672B6000C86824192C44FAD8EDF068C6DA",
            INIT_RAM_36 => X"28142339BCE66FB75A883822110A8665B4BB6D170181B0926BC1C990726A3C94C160422C",
            INIT_RAM_37 => X"0E0907A3533198CC9D6EC7AAD56ABC7A9F379B994383D33198CC66000000000000000050",
            INIT_RAM_38 => X"4A00299D6B726C3612E8D4B43E0F0470CAC65B294295BCDC8BC75BADA74A81C122753A24",
            INIT_RAM_39 => X"8CA62A1202806828140A04C3612092CFAD1CF2F97CBE5F2F57AB54DDEEDB4592DA58CC66",
            INIT_RAM_3A => X"00000000000000000000160A0584C466A7D3EA772B551D0E8733996D07046120DC66B298",
            INIT_RAM_3B => X"59A513A1C0E155BB1E4E954CC6633198CC9673399BD1EABC7A3CDD4E3992C6E4B198CC66",
            INIT_RAM_3C => X"F1EECB01B2A870381C2AA5401DEB7270361BACF27C1E0F0745AA65632D8391B95E6B35E3",
            INIT_RAM_3D => X"12030480C0D964B258282633258090B028140D85024120975BCBE5F2F97CBE5F2D566919",
            INIT_RAM_3E => X"4B259BCDE6EB79BC9400000000000000000014285B2C848160B05854B66455ACDE4AB319",
            INIT_RAM_3F => X"5B2D86A5CF1C8AB5E399870B8BE12070383D6EB78DC6633198CC66331B92C9632994DC96"
        )
        port map (
            DO => promx9_inst_12_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_9,
            RESET => reset,
            AD => promx9_inst_12_AD_i
        );

    promx9_inst_13: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F2F97CBE5A6064339BF1F8C001C1186C24120E154874CCF2B0361A6D783C1E0F0686261C",
            INIT_RAM_01 => X"2C160B05028141A29B0603018430D86C60582C46530301605028140D86C245AEB797CBE5",
            INIT_RAM_02 => X"33198CC6633198CC6633198DC663297048950000000000000000000016542DA8CB44B058",
            INIT_RAM_03 => X"6D747C1E0E8F4F446532AD94A13DDD6F37196D830385C6EA50CC552A995BCDD4B198CC66",
            INIT_RAM_04 => X"0D86CB59EF2F97CBE5F2F97394C10A6D35E4ED66850230D84824120D8D52C9AEB3103612",
            INIT_RAM_05 => X"00000000070C6A3319640C0A09828241B40C0E030381B0D8A050502C340601B2D86C2814",
            INIT_RAM_06 => X"33198DC966F378DC6633198CC6633198CC6633198CC552A998CC66000000000000000000",
            INIT_RAM_07 => X"090712C5AEB290241B8CEC3C1E0F07273CDC0A2956C148DF8E459B8C9506A1C12275BA1C",
            INIT_RAM_08 => X"2C140B25A0905028140916FADDEF2F97CBE5CE679B6192D26AB7E3F1C68421B0906C381C",
            INIT_RAM_09 => X"0000000000000000000000000282814232E168B8632C848464A8542183046230C8A0A028",
            INIT_RAM_0A => X"A8C683835331553ADE32998CC66372763C9D37198CC6633198CC6633198CC6633198CC66",
            INIT_RAM_0B => X"ED468421B0D8F4381C2188CCC5AF3B70241A8CF47C1E0E8E8BAD13099958C355278F951A",
            INIT_RAM_0C => X"06070A8542D168005814140322816050281B0906CB59CF2F97CB9C9A16432598DD6FCDE3",
            INIT_RAM_0D => X"33198CC6633198CC6600000000000000000000000000000285C31A70B85C2A16CC65B49A",
            INIT_RAM_0E => X"2D8718C650DF53A751ACD65C6940E0D4CC958F2F8CA6633198DCDE8F2F92C6633198CC66",
            INIT_RAM_0F => X"2D04833A56D793D9E3ED464501B0D98C4223060706A1ADF474321A6D783A3E0F076F391C",
            INIT_RAM_10 => X"8CC6632C88CC6632430E07038430E0A0502800160B05A0A05036120904A99E5EB44F1C5A",
            INIT_RAM_11 => X"37259BCDE4B1B8CC6633198CC6633198CC350000000000000000000000000000000000A1",
            INIT_RAM_12 => X"50F4BA5E0F0727ABE709050CA650A54F23AAACE6644BB2A1547A352AAF9BC9637198CC66",
            INIT_RAM_13 => X"0DB73AD9C2D36CB2192C965C753CE793DBE3F1C683212DB6D8460C0E070CC5ADF454421A",
            INIT_RAM_14 => X"0000000000000000000046633198CC65B40C2A0E8A8430D00000002C16042140A0503623",
            INIT_RAM_15 => X"33198DCDE6F1B8CC6633198DC966EAF9BC9633198CC66330D4381C000000000000000000",
            INIT_RAM_16 => X"06070CC9ADF16C321A2D78FC1D2F07833DE72D86C6A650A273A9C9E4C65769473198CC66",
            INIT_RAM_17 => X"2C14026140A05028142E6F9B4190C96C2459CCAA7D8DAF37B3D9E3F1D64501ADB2F4180C",
            INIT_RAM_18 => X"0000000000000000000000000000000000002CC6633198CC6536544D2CD349B000000000",
            INIT_RAM_19 => X"F06C1B49D21A58CC6633198CC664EC792C6633198CC66332592CDE8F378CA3D06070381C",
            INIT_RAM_1A => X"F1E68421ADB070180C060D52CB3B729042210CF73A5E3F078337E78A848289D0A073B9D2",
            INIT_RAM_1B => X"6D36976000000000281400058140A05028126E16032190C864B399A846FD934F67B3D9E3",
            INIT_RAM_1C => X"2E275BADD6EB752C3D0000000000000000000000000000000000004C46633198CB8536D9",
            INIT_RAM_1D => X"F384836650A17227E3E978332BB4A96D2C6633198CC66331B9BADE4B198CC662A9547A5C",
            INIT_RAM_1E => X"887B3DB5BF27B7D9E4F1F8CB01A32830180C0E154C71DB7270321910D6BA5E3E8E8BB7E7",
            INIT_RAM_1F => X"2CB2232E18CC6632D98CC6542000000000000016828140A0B032592C80032192C96793D1",
            INIT_RAM_20 => X"6EB74DC6633198CC6633198DC6E6EB76BB5D000000000000000000000000000000000000",
            INIT_RAM_21 => X"10B87B7E3E974F45E7F396C36350A273B9E3D0F83C1A12DA54469533198CC6633198CC6E",
            INIT_RAM_22 => X"0006432D92CE67C1E0A9F93DB9CF6E6BD9E3F1F8DB41A1D0F4AA351EA5843BEB7358341A",
            INIT_RAM_23 => X"00000000000000000000469A31A68C6633198CC645000000000000000502814118640028",
            INIT_RAM_24 => X"2E2597A9533198CC664B259BCDD37198CC664B2557AB399E6FA7D3000000000000000000",
            INIT_RAM_25 => X"33251B96E9349832194D386B5E3F1E8739E7F3B7024142E173C7E3F1F83C1E0AD1512A94",
            INIT_RAM_26 => X"0C850285C00000000000086B298D0F83C1E0EA7B3DBE4F1F2BD9ECF1E6FD80009194CC66",
            INIT_RAM_27 => X"00000000000000000000000000000000000050A44A0918CB85B2A18CB852200000000000",
            INIT_RAM_28 => X"F1F4BC1E0E8CD0CA5C4A8E92B3C9E2F52C96332552B1EAEB767933CE66FC7E3F1F8FC7E3",
            INIT_RAM_29 => X"F1F8FD91A1406D2C664B086DD6E63395761970B6633DBF1E87CF9EF3D1824144E2CFB9E3",
            INIT_RAM_2A => X"8CB85C2000000000004D050360000000B00000442A199E8F83C1C9CDFB3D9ECE572BC9EC",
            INIT_RAM_2B => X"AE66FC7E3F1F8FC7DA0000000000000000000000000000000000000000122904C3852151",
            INIT_RAM_2C => X"F3F9C24130DD33B9E3F1F8FA3E0E8E65669612258B85B9E572B7335EAF57ABD9E4D3A99C",
            INIT_RAM_2D => X"D57B3D9EDD4727DBECF278F77ED488A024632D49ADD6E6339656596CC663392F1F73399E",
            INIT_RAM_2E => X"00000B29A2C1A1B2988CC65420000000B1992D96D30910000000002CF4733E0F0783C192",
            INIT_RAM_2F => X"F1F8FC79BCDEEF37D4EA74FA7DAF1F8FC7E3000000000000000000000000000000000000",
            INIT_RAM_30 => X"4CC663319EDF9739E7F3F9E381B09E6FC7E3F1F8FC7D1F0666689D33150A8962A16E79E4",
            INIT_RAM_31 => X"ACF83C1E0F0747C1C9E9F53D9E4E8763DB9CF666FDBEDCE160005B6B5BADD6E6B476B6DA",
            INIT_RAM_32 => X"00000000000000000000000B0001426531198CC64B000000A2B3D159D663200000000000",
            INIT_RAM_33 => X"2A9B8DC2432A58B69A6DE6F37E3F1F8FB5E3ED74FA7D4E9F6BB5E3000000000000000000",
            INIT_RAM_34 => X"6349ADD6E93577375C70C66331ACD78FADE7F3F9FCE120A2CFC7E3F1F8FC7E3E978234BD",
            INIT_RAM_35 => X"905640000488000058ACE87C1E0F0783C1E0F26ABD9DAE8743DB5BF6FB339A4F346948C6",
            INIT_RAM_36 => X"0000000000000000000000000000000000000000000001416120E170B84B02800162A3E0",
            INIT_RAM_37 => X"F1F8FC7E3D174BA31A4B1B9CC964A891BD1E9E36E575BCDF8FC7E3F1F8FA7D3E9F53A7E3",
            INIT_RAM_38 => X"6DFB739E6D2FB5CAC6632DA4D6E72F77D99BADC663392AD78FBDE7F3F9FCEA40D84BB9E3",
            INIT_RAM_39 => X"8CA41420000367C1E0D0801315A2C16122008CF47C1E0F0747C1E0D56A7D9CAEC74377DD",
            INIT_RAM_3A => X"ED78FC7E3E9F4FA7D400000000000000000000000000000000000000000000028001B2E1",
            INIT_RAM_3B => X"F3F9E8D8E0906E27E3F1F8FC7E3F1F4BC1E0A9B98ED565F2F8B89CAEE7B379BCDF8FC7E3",
            INIT_RAM_3C => X"D5727DBCAEC763B55C5DFB7CDEDF6F9A367E32B19AD6E8AFB7DBE4F23863392C978FBDE7",
            INIT_RAM_3D => X"000000000000A120E18CC6800004C747C1C92C44332582C46450A1E8F83C1D1F0683C1E0",
            INIT_RAM_3E => X"4E2B2BB9ECE673B5E3F1F8FC7E3F1F8FB5DA000000000000000000000000000000000000",
            INIT_RAM_3F => X"F6C663392D1773B9E7F3F9F3C122D848259BA9F73A5E3F1F8FA5A0CCD6ABCCE9B5BA6CBE"
        )
        port map (
            DO => promx9_inst_13_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_11,
            RESET => reset,
            AD => promx9_inst_13_AD_i
        );

    promx9_inst_14: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"F078393E0D8747C1D1F0543BBCAE874394BB6DE93CDE6F36DBDA24261954AD68EFB3C9EC",
            INIT_RAM_01 => X"0000000000000000000000000000000050D970B212200ACF83C0E08CE64B0988C96535B0",
            INIT_RAM_02 => X"D0ED2A75DB74FADD6E9F5799CDC6E5773D95CEE73A7D4E9F4FC7E3000000000000000000",
            INIT_RAM_03 => X"12050CAB6AEFB3D9ECF266E335AF1F8FC7DEF3F9D9C9C0D8482412CE36BA5D2F1F4BC7DB",
            INIT_RAM_04 => X"D0AA633222D26B33E0D0D43C1B08878341A0E896A37CAE8743532B6218FCDA5F3696781C",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000598CB8400A9F07834159",
            INIT_RAM_06 => X"4D44E99A1E974BA5E3F1D6B7D6EB75BADD6EB75BADD6ECF475B8DCAED772B9CDA673A7D4",
            INIT_RAM_07 => X"4D16BCDB6ADED8B6541205038B6D2F77D9ECF266E3392F1F8FCB9CF3F9EDC6E0D86C2412",
            INIT_RAM_08 => X"70A6001A1F074733E0ACE6534126D687A3507068342E0E8E8221C954848259BD4F43A522",
            INIT_RAM_09 => X"8EC55B91BA9CD2BB9C000000000000000000000000000000000000000000000000000090",
            INIT_RAM_0A => X"EB79FCEDE3290C46120D9693553D0F47A5E0E978F358EB75BADD8EB75BADD6EB763B3D9E",
            INIT_RAM_0B => X"2D06C24A1EC74BB9910D86AB812626D8460C261302865AE793D9ECF6791C392F1F8FB9D6",
            INIT_RAM_0C => X"00000000000000005070800B1D1F0686A5516D17036DACCD41C0E0D8681C15088382A098",
            INIT_RAM_0D => X"B75BADD6EB75BADD6EB75BB1D9EAECD2375B000000000000000000000000000000000000",
            INIT_RAM_0E => X"F67B1C392F1F8FC7DEF3F9EDD3E3708D2C1209048241289F27A351D0E87A5E3C763ADD6E",
            INIT_RAM_0F => X"88381C0E0883813012090482412D4F73C7920D26D881A31968360C0E050281C9A793D9EC",
            INIT_RAM_10 => X"0000000000000000000000000000000000002C8A241D16C97166140A06CB45A68381C150",
            INIT_RAM_11 => X"A654AA552A9556DD6EB75BADD6EC75BADD6EB75BADD6ECF67B3D9E000000000000000000",
            INIT_RAM_12 => X"0E0B028142E79BD9ECF27B6335AF1F8FC79CF3F9FCEBE6F1B898650906C241B0916AB59B",
            INIT_RAM_13 => X"0D84824A14C38220E0703822110702A424120906C245AD4F4BC7DB34B8CB41B09048360C",
            INIT_RAM_14 => X"0000000000000000000000000000000000000000000000000000282C0A332910A0502814",
            INIT_RAM_15 => X"21848241209048B2DA8E3558CD59363ADD6EB75BADD6EB75BADD6EB75BADD8ECEE773B9C",
            INIT_RAM_16 => X"4D36DC6120D86C461C0E13028140A2B3C9E4CE571C319F1F8FC7DBF2F9FCF3E6F1B93A66",
            INIT_RAM_17 => X"0C801A05B0E050281409069229850B81C0E070381C0E05484824120904824DCF1F4BC7E3",
            INIT_RAM_18 => X"B75BADD9EC76773B9D000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"AA557CFBE3B258CC6E3310C24120908C24124D2CE2AB65B2964D6EB75BADD6EB75BB1D6E",
            INIT_RAM_1A => X"09048294CF1F8FC7E3A9D0EA65B0908C461C1E89028140A06F39ECF3369C2E1EDF8EA953",
            INIT_RAM_1B => X"00000000000000000014001202C0A050281B09164B45A54B81C0E088381C0A909048241B",
            INIT_RAM_1C => X"935BADD6EB75BADD6EB75BADD6EB75BADD9E000000000000000000000000000000000000",
            INIT_RAM_1D => X"8DB11B5198D772A8DC4E5522B1D6F198CC6633258461209048241209048B4B4632D96CD5",
            INIT_RAM_1E => X"7038152120904824120906C29E3F1F8FC7E3F1A6FB8C40D890380C0E19898140A051B91B",
            INIT_RAM_1F => X"0000000000000000000000000000000000000016120140A050281209068365970285C0E0",
            INIT_RAM_20 => X"0906DCA9C4EAD98CB66331A4D6EB75BADD6EB75BADD6EB75BB7DBE000000000000000000",
            INIT_RAM_21 => X"060D4CC4C0A050B85B2D37024DA9864BB65B6216D88DD26198CC66331992C4C090482412",
            INIT_RAM_22 => X"59A74A8982D245C1507036824120904824120A05239E3F1F8FC7E3EE48BC6941188C180C",
            INIT_RAM_23 => X"000000000000000000000000000000000000000000000000000000000A0B4430D050281B",
            INIT_RAM_24 => X"33198CC663288C24120D84826B65B2D96CB66349ADD26B75BADDBECF67ADD8EB763AA954",
            INIT_RAM_25 => X"F1F73C6240606C183D0E030CC661605058120916C245A8CB8335532A0F4B8244E954CC66",
            INIT_RAM_26 => X"000A1325A2E0502812CF194B4122CB8241207017024120D86C24140A073B9E3F1F8FC7E3",
            INIT_RAM_27 => X"A9E6F699DCEE773BB4000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"50830381C0E070CC6633198CC6633258CA230904824125B3196CB65B2D96D26B75BADD54",
            INIT_RAM_29 => X"0A273C7E3F1F8FC7E3F1F8FB61C0608C183506070CC66330B0585B2D048B4122CB41C19B",
            INIT_RAM_2A => X"0000000000000000000000120591186C365BDA08C365A88383A0E06E048B812090483614",
            INIT_RAM_2B => X"5B2D96CB65B3564D6ECF552B3A9E86A351A8000000000000000000000000000000000000",
            INIT_RAM_2C => X"6D0483612092A5C0E0AD268380C0E0306A6633198CC6633198CC9526130361209171ACB6",
            INIT_RAM_2D => X"4E170B6120904828140A2D3CBE3F1F8FC7E3F1F8EA80C06070181C330306A66331B8584C",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000050682E050371C6687086D0ACEA750E0",
            INIT_RAM_2F => X"3286846120D84CB8D65B3196CB65B2D98CB6935BB3D9DC9567A1D0000000000000000000",
            INIT_RAM_30 => X"2A9987A663319898768D46424120904930E070260B81C0E030386633198CC6633198CC66",
            INIT_RAM_31 => X"1210CB3A09074352B32DA7424120D86C28650A533BDE3F1F8FC7E3F1F8DB80C06030180C",
            INIT_RAM_32 => X"00000000000000000000000000000000000000000000000000000000000009A1197025BE",
            INIT_RAM_33 => X"33198CC6633198CC6633258862421AB0B8134E3196CB65B2D96CB65B2D96CD5B767B69AA",
            INIT_RAM_34 => X"F1F49380C0603038351E998AA6633198CC656DF41B4592C968B4E088441423D2D830183D",
            INIT_RAM_35 => X"0000000282D849B915060EAB3D8D474240D62E35424120A06CCA650A557BDE3EE78FC7E3",
            INIT_RAM_36 => X"5B2D96CB652AD9AB15000000000000000000000000000000000000000000000000000000",
            INIT_RAM_37 => X"70381C05A1D16C180C2A998CC6633198CC66331992C630E09098D652A956CB65B2D96CB6",
            INIT_RAM_38 => X"0A67BCFDCF2F8FC7E3E9749380C0E030183D0E1997A66332F4CC665EF43B0D12CAA424E0",
            INIT_RAM_39 => X"0000000000000000000000000590904B1C240636F41D8E874240D64E97024120A1716C65",
            INIT_RAM_3A => X"4EAD96CB65B2D96CB65B2D96CB65B319B922000000000000000000000000000000000000",
            INIT_RAM_3B => X"4B68393A154B81525970381C0D05D964B81C0E1B8CC9633198CC661A8D4CC66260303824",
            INIT_RAM_3C => X"5299436121A9956CA509DBBCFDCF2F8FCBE3E9782865B06030181C332F666662AACD2C95",
            INIT_RAM_3D => X"000000000000000000000000000000000000000000019092CE2A0C0E683B1D0E8742B4B6",
            INIT_RAM_3E => X"33154383533090181C262756CB65B2D96CB65B2D96CB65B2D96CD5000000000000000000",
            INIT_RAM_3F => X"1AAF6B2B35EA59B6955EE8795A0CD381C05970565C1194C269305B0E0F5BADD6EA54CC66"
        )
        port map (
            DO => promx9_inst_14_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_13,
            RESET => reset,
            AD => promx9_inst_14_AD_i
        );

    promx9_inst_15: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"4DF6393D0E864626B65B194B81B32A956CB609F9FCFE5F2F73CBDCCCF83931A06030380C",
            INIT_RAM_01 => X"00000000000000000000000000000000000000000000000000000000000000000638480C",
            INIT_RAM_02 => X"8D8912934DA551BA6E33198CC0C0E0D4181C121D93AA55B2D96CB65B2D96CB65B2D96CC6",
            INIT_RAM_03 => X"AD727C1D12D830869B0E25AB3594A2F6B2966DE6741E3E4D69C0E054B82A7198D381C0E0",
            INIT_RAM_04 => X"0000000004D4D0180CACF4393D8E8566A6B65B294B45C52B198C6509F9FCFE7F2F8FABDC",
            INIT_RAM_05 => X"5B2D96CB65B2D96CB6000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"703833919CE481C0E07046A691BCDF8FC7546EA54CC662A870180C06070987E5B2D96CB6",
            INIT_RAM_07 => X"32DBBCFE7F2F8FCBE58CF8361E08D10CA8D94D10EB7D099B6F3533ACE6793CAED78DC110",
            INIT_RAM_08 => X"000000000000000000000000000CF170180CD0F4393CAEC54EA6B65B318269C52AD98C23",
            INIT_RAM_09 => X"0E030181C261F94AB65B2D96CC65B2D96CB6000000000000000000000000000000000000",
            INIT_RAM_0A => X"ADF6393C9F1F8FA6E08D38233E6CE7B1B3108846A2152CE78FC7E3EE551BA95331986A0C",
            INIT_RAM_0B => X"632D8B8D632AD98C1216457CFE7F3F8FCB9E8D56661E0AC86966DA8CC6741D8CD56667A0",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000B38A870180CADEA393CAE856626C6",
            INIT_RAM_0D => X"F1F8FB9546EA592C6606070180C0E070987E6B2D96CB65B2D98CB6000000000000000000",
            INIT_RAM_0E => X"8CC6741D0D4726B5A0D0743A1DAED76BB55968671319BF6793DB1A70347BBD3EDF8FC7E3",
            INIT_RAM_0F => X"99F6B95A1F1EA22AB65B2D98C65632D98C1221B77CFE7F3F8FCBE7A94C191A9A816932DA",
            INIT_RAM_10 => X"00000000000000000000000000000000000000000000000000000000000019D12030181C",
            INIT_RAM_11 => X"F256A33B4EDF8FC7E3F1F8FC7E3F1E6E87345E9987A1C0E0301824261F96CC65B2D96CB6",
            INIT_RAM_12 => X"EAA4260C8A81A0A1198CC6633D8EC76341D8EC763B1C9F1F8FC7E388467DB1AEA7B3D9EC",
            INIT_RAM_13 => X"0000166DD06030381C59F8F93E3E576AB4D5633196CC663319AC430D49B7DE7F3F97CB9E",
            INIT_RAM_14 => X"0E070484C3F2D96CB6000000000000000000000000000000000000000000000000000000",
            INIT_RAM_15 => X"E9B8235EDF27B3C9ECF27B3DBECEA753C7E3F1F8FC7E3F1F8FB99AAD46AA6DB6E970A854",
            INIT_RAM_16 => X"4ECDF3DE7F3F7BB9558DA6130986C940B0908CC663351EC763B1D8EC727A1D0F1F8FC7E3",
            INIT_RAM_17 => X"000000000000000000000027C240E031661C59CCFC7E3ED78F951C633196CB65B2D98C12",
            INIT_RAM_18 => X"F1F8F45A0D0E6733598D2EC863D2A130987E000000000000000000000000000000000000",
            INIT_RAM_19 => X"EC68393D0E578FC7DAF1F4DC153F67B3D9ECF67B3D9ECF6777A9DBF1F8FC7E3F1F8FC7E3",
            INIT_RAM_1A => X"9A3196CB65B2D98C1A9339AAFE7F3F9F39553426140A048160B030645463319D476393D8",
            INIT_RAM_1B => X"00000000000000000000000000000000000000471880C06072B60CD22CFA7D3F1F6BC7D3",
            INIT_RAM_1C => X"E9F8FC7E3E978FC7E3F1F8FC7E3E9747C1E0E8E8733594D18CB623000000000000000000",
            INIT_RAM_1D => X"4838633198CEA393DAE872B95C9EC78FC7E3F1F6B34E0CDF93D9ECF67B3D9ECF6793A9D4",
            INIT_RAM_1E => X"6DCCE679DE9F4FA7D3CDD516CB65B2D98C236EC9A6FBEF3F9FBD554C28130984C160B0E1",
            INIT_RAM_1F => X"00000000000000000000000000000000000000000000000000000000678380C0603336B3",
            INIT_RAM_20 => X"F6793D9ECF67B3C9D4EA753B9E3EDE87C7E3E978FC7E3F1F8FB7A1E8F83C1E0E8E86B2DA",
            INIT_RAM_21 => X"4C26130984C160B0C88CC663319CD567A1E3E5727C7DAE4F8FC7E3F1F8FC7CA7066FDBEC",
            INIT_RAM_22 => X"A62B0180C06032679B59EEDB79CDF74F2BD3AEF4E2AC65B2D98C5C21D3E9EDDF3F9FCF9E",
            INIT_RAM_23 => X"E974BA5D1E8F83C1D1000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"F1F8FC7E3CD382A7ECF67B3D9ECF67B3D9E4EEF53A7DBF1F8FA3D2F1E8BA3D2F1F8F45D2",
            INIT_RAM_25 => X"0DD3CB61CF3F9FCFE734260D0685096060908CC6633198CF6B35C9F1F2BB5E3F1F8FC7E3",
            INIT_RAM_26 => X"000000000000000000DF070180C0E08E67E399E6F772BDA6D355BEAA552A6D5632D96C5C",
            INIT_RAM_27 => X"E8F4BA5D1E8F47A5D2E8F47C1D1E8F47C1E0000000000000000000000000000000000000",
            INIT_RAM_28 => X"F1F8FB5E3F1F8FC7E3F1F8FB5E3F1EEDB35AF6FB3D9ECF6793D9ECF6793D9D4E9F73A5D1",
            INIT_RAM_29 => X"DF5523B345B3196CB60916C481C8AF9FCFE72C260B09048161325870C6633198CD67C7BB",
            INIT_RAM_2A => X"00000000000000000000000000000000011C8A90C180C0615135E3F1F6BB59BCDF9F69B4",
            INIT_RAM_2B => X"F67B3D9ECF2753A9D3E9783C1C9E8F83A3E0E8F83C1D1E8F4743A1000000000000000000",
            INIT_RAM_2C => X"6446632DA8CCAEA3E3F1F8FB5E3F1F6BC7DAF1F8FC7DAF278FC95368777C9E4F6777D9EC",
            INIT_RAM_2D => X"ED78FB5D4E9ED3CFB4DF7562B556AAD93AB621848489611F9FCFE750960B0682C1A0B0DA",
            INIT_RAM_2E => X"0000000000000000000000000000000000000000000000000001D60D870181C06071355B",
            INIT_RAM_2F => X"F646AB7E4F67B3D9ECF67B3D9ECF67B3D9DDF275355C9CCE87A3A1D0D4AA552A65322B15",
            INIT_RAM_30 => X"6D140B0582C160609B8CC6632DA6D3677759F1D6FC7E3F1F8FC7E3F1F8FC7DAF1FB337EC",
            INIT_RAM_31 => X"11830180C2A10D6719F1F8FC7B4DA74F69E7CE79F3CC672AD99CB62E049CCE60E5BBCFE7",
            INIT_RAM_32 => X"EA6573B1D6AAD96CB600000000000000000000000000000000000000000000000001674C",
            INIT_RAM_33 => X"F1F8FC7E3F1FB3D9ECF6777C99BF27B3D9ECF6793D9ECF67B3D9ECF2777C9ECEEF77C9DD",
            INIT_RAM_34 => X"4E84A9E3D06133CF6E8D960B030280C0B0124D46633195DB69B5BBF1B6E67E3F1F8FC7E3",
            INIT_RAM_35 => X"0000000000006698DC1D03136544D1513522ACE6BC7D3F3EFBA9D5F3E7BCF556AAD93A7E",
            INIT_RAM_36 => X"EEE76BB5DCAD773B5DB7455AAC6632D96CB6000000000000000000000000000000000000",
            INIT_RAM_37 => X"99CCCA933DDF8FC7DAF1F8FC7E3ED78FD9ECF67B3D9ECF27B3D9ECF67B3D9ECF27B3D9EC",
            INIT_RAM_38 => X"F3F9FCFE7A32D96CBE5B3352C1C060733D266E260B04318168B0214AB6632DA6CA6C869B",
            INIT_RAM_39 => X"00000000000000000000000000000087BC9B0D90E449BD026D36D98CF8EA3E3DA79FCF9E",
            INIT_RAM_3A => X"F6793C9DDF67B3D9ECF27772B3472B55AAC652B558CA5632D96CB6000000000000000000",
            INIT_RAM_3B => X"1D071349B4DA69365421CCE663D59D6FC7E3F1F8FC7E3F1F6BC9ECF67B3D9ECF67B3D9EC",
            INIT_RAM_3C => X"8CD6AB551F1E73CFE7F3F9FCFE7F3C556C9D37274380C06031BB6E6E160A023218E8B458",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000C96FCA9B0DACEB359CCE81B4DA",
            INIT_RAM_3E => X"F67B3D9ECF67B3BBECF67B3D9ECF67B3D9DDF67B3C9ECEEE563B1572B19AAD5632D96CB6",
            INIT_RAM_3F => X"5F160602C06150183A10950A89B1D070861C06070A8540615167BBF1F8FC7DAF1F8FB5EC"
        )
        port map (
            DO => promx9_inst_15_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_15,
            RESET => reset,
            AD => promx9_inst_15_AD_i
        );

    promx9_inst_16: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"12AA9C0DCB0154AAA2B032E471D8EC88970381C0E070381C0E8802140A346F49C4E17153",
            INIT_RAM_01 => X"5528DB6D98580804020000000000000000000000000000000000000000000006532D149C",
            INIT_RAM_02 => X"75DBCD46A351A8D46AB85C25B7096CB6E17096CB6E170B80B25B70B85C2E170B85C0E42C",
            INIT_RAM_03 => X"048D465389C1ECF66B5D22E24D19C4E270F41B3AA70F4596C271389C4E1E8F49C4E271B0",
            INIT_RAM_04 => X"00000014A0041E0EEAB1BADC09D2AB7128C98A34EACDB0AB91284B25C1A070381C0E1544",
            INIT_RAM_05 => X"B85C2E170968B1469345A4E1744018080402000000000000000000000000000000000000",
            INIT_RAM_06 => X"9C4E360367A4E271389C6C2E06A351A8D5A996DC2E170B85C2E170B85C2E12DB85C2E170",
            INIT_RAM_07 => X"45C2A070381C0E070301958F67B3D9ECF67BD1B5218CB7A4E271389C4E271389C3D27138",
            INIT_RAM_08 => X"00000000000000000000000000062B159625B1B8DC0E0253248844A8C51169B69B5536CB",
            INIT_RAM_09 => X"B85C2472371B8DC6AB96DC2E170B85C058A3A20080402010080402000000000000000000",
            INIT_RAM_0A => X"9C4E270F49C4E271387A4E1C6E3594E270F47A0D9D6EB351AA5A6A71DBEE170B85C2E12D",
            INIT_RAM_0B => X"A2449968B8580DA6CB85C1D888425A120703834282A353D9ECF67B68B4E24D1564E270F4",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000006292E3563B1B8DC0E064D121544",
            INIT_RAM_0D => X"B84B65B2D96DC2E02CB84B4E52DEBA2B07832272993D771CB6E02C1642A1543048240602",
            INIT_RAM_0E => X"65B1A94D1ED3D271389C3D271389C4E271389C4E1E8944A2AB61389C3D1647475BAB532D",
            INIT_RAM_0F => X"12B8DC0E02AC2A8944A21299602658281506A2312894445313910A81F4C2A283D9ECF7DA",
            INIT_RAM_10 => X"1628E0AC6633198C8A000000000000000000000000000000000000000000000A54292763",
            INIT_RAM_11 => X"75CE270B2B91CAE16FB85C2E17096B8DC6E371B8DC6E3719C9C784C1E0F0644C1F2A24E3",
            INIT_RAM_12 => X"25429B228141EDA2CB6582694CB68E8D59387A4E271389C3D271389C4E270AA2272928E3",
            INIT_RAM_13 => X"0000000C500316AD63B1D81C0E064B168944A251390026500C0602013128944222290A85",
            INIT_RAM_14 => X"42E0F0783C1E0F068569BC9B8CB65B2D96CB000000000000000000000000000000000000",
            INIT_RAM_15 => X"9C4E1E8F43291306444544DD6F45526DC6E371CB647D771F5F0983C1E0F0783E5227AEE3",
            INIT_RAM_16 => X"A211289442221615CA6232D26E43468D8C0904C2994CA68B2DD4F495BA959387A2B154F4",
            INIT_RAM_17 => X"000000000000000000000000000A532F929C12D813AE0895128944A211188C4015100402",
            INIT_RAM_18 => X"C1E0F0783C191088448960F0783C1E0F078342E19C8CB65B2D96CB000000000000000000",
            INIT_RAM_19 => X"7638E2738D42C9C665594E0CAAA591951583C1E0D14E3592288844221130912C1F5FAF83",
            INIT_RAM_1A => X"A251188C40100805446251288C5C1E0D0B0A65A168685ED76914854280A1586A1B2F46DB",
            INIT_RAM_1B => X"0000000000000000000000000000000000000000000000022E156312D8DC0E04EB268944",
            INIT_RAM_1C => X"C1E0F0783C1E0CAB83C1E0F0985452151244C22148844C19110A4422619991365B2D96CB",
            INIT_RAM_1D => X"A182804CA012298CD3A500219199C465D6948A2A9D71389C4D2889C1E0C89834DA6F0783",
            INIT_RAM_1E => X"B1D8EC09D4EB711344A25118B440100804C5A25118A44C1A16149342C28040AA1B181202",
            INIT_RAM_1F => X"42E0E16CB65B2D96CB00000000000000000000000000000000000000000000062921149C",
            INIT_RAM_20 => X"C1E0F07832244F07832260F0783C1E0C8844C1E0C894A0030D89894522E88852260D0ACB",
            INIT_RAM_21 => X"A9C16170601A49940A0142A88020180D14CCA500000006538E94DB89A2A2713C21130783",
            INIT_RAM_22 => X"0000000006533114D1B1D8E45606E75C9544A25108944A1A159744A2317078342C2B0CCB",
            INIT_RAM_23 => X"003119686A2227068524214890565B2D96CB000000000000000000000000000000000000",
            INIT_RAM_24 => X"003111544449130783C1E0F0783C1E0F0783C1E0F0644C1913078342F288844A20000000",
            INIT_RAM_25 => X"62E0F06C58532D268B62B4C00D36532C00CA048249002010299856628000000000029400",
            INIT_RAM_26 => X"0000000000000000000000000006552A15C9B1D8EC722B035596CB83B2E0D0582B2E8844",
            INIT_RAM_27 => X"E530F0A894532D86000000000C369B111583659210ACB65B2D96CB000000000000000000",
            INIT_RAM_28 => X"4A31400000000000000000296C6C4F291783C1E0F0644C19130783C1E0F0783C19111383",
            INIT_RAM_29 => X"82B2D96CB65D118A85C1E0D8BD66180000C5A5328000045A4C00002442C010B013312800",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000C500344908A69D8C4A259136D98CB",
            INIT_RAM_2B => X"C1E0F0783C1A2588852262400006230996C300000000000319868A22331958665B2D96CB",
            INIT_RAM_2C => X"0025194C5053298CD30000000000000000000000000C30022587CAC1E0F0783C1E0F0783",
            INIT_RAM_2D => X"EA251A8D369B4D24C66332D97058312216CB42C2996000000000000000000000022D8A00",
            INIT_RAM_2E => X"42D118AD385B2D96CB000000000000000000000000000000000000000000000A50010ACB",
            INIT_RAM_2F => X"2260F0783C1E0F0783C1E0C8983C1E0D88C4451129400000000000000000000000000000",
            INIT_RAM_30 => X"000000000000000000005298C006322D8A00000000000000000000000000000005298886",
            INIT_RAM_31 => X"00000000000001954A65A2DA8DA6D351168B45A2E0D068332A168BEB32C0000000000000",
            INIT_RAM_32 => X"00000000000000000061A2C000062A4996CB000000000000000000000000000000000000",
            INIT_RAM_33 => X"00000000000002960045E0F0783C1E0F07832260F0783C1E0F120061E251589000000000",
            INIT_RAM_34 => X"00000000000000000000000000000000000000000000000001A600000000000000000000",
            INIT_RAM_35 => X"00000000000000000000000000000000014A003158B86C312090CB65B2D969365B2E16C6",
            INIT_RAM_36 => X"0000000CB65A3000000000000000000000000030C0000000010A92000000000000000000",
            INIT_RAM_37 => X"0000000000000000000000000000000186006260D16442260F078344E0F0644C1E0D12C3",
            INIT_RAM_38 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"0000000000000000000000000000000000000000000000000000CA003280000000000000",
            INIT_RAM_3A => X"C2227078442E0F0789000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"000000000000000000000000000000000000000000000000000000A522584C9C4E0F0644",
            INIT_RAM_3C => X"A50000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"00511848B61A28888A42E270783C4A170644618000000000000000000000000000000000",
            INIT_RAM_3F => X"000000000000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => promx9_inst_16_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_17,
            RESET => reset,
            AD => promx9_inst_16_AD_i
        );

    promx9_inst_17: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 9,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"0DA6FB1A8D06A753226CC7337198CD673DE7F3F9FCFE7F3F9DAAB63B1D8981C061546B6E",
            INIT_RAM_01 => X"D2E573B3E72AD96CB600000000000000000000000000000000000000000000010B73AC1A",
            INIT_RAM_02 => X"6DEEFC7E3F1F8FC7E3F67B3C9ECF2793D9ECF2793D9ECF6777C9ECF67B3D9ECF67B3DBDD",
            INIT_RAM_03 => X"5B1B92C0C2A998CCDE4B164602C06030181C1E88C181C2A10C180C06030381C060301843",
            INIT_RAM_04 => X"0000000280053298230936FB1D0D4EA3A9D28CB6E68E1A1D6E359ECF67BCFE7F3F9FCED5",
            INIT_RAM_05 => X"F67B3D9ECF27772B1D8AC75CAD5632D96CB6000000000000000000000000000000000000",
            INIT_RAM_06 => X"06030863D0E030180C0610E67E3F1F8FC7DAF27B3D9ECF67B3D9ECF67B3D9E4F67B3D9EC",
            INIT_RAM_07 => X"8AF57CFE7F3F9FCFE763338CC6633198CC6626268A0140E030180C06030180C06070180C",
            INIT_RAM_08 => X"0000000000000000000000000000CD56381B0926BB1D8EE74BA3DCE9B464D1A6DB6A351C",
            INIT_RAM_09 => X"F67B3379BE9F4FA99CF27B3D9ECF67B3BB956AAD96CB65B2D96CB6000000000000000000",
            INIT_RAM_0A => X"06030181C06030180C0E030C6DA2A030181C0E0F528DBF1F8FC9E3E9EEFD9ECF67B3D9E4",
            INIT_RAM_0B => X"F1E49B9156D319B6DC72D3339DECF77BCFE7CF274FC6E33198CC6616068602C12030181C",
            INIT_RAM_0C => X"0000000000000000000000000000000000000000000000CE79C6120926BB1D8E978FB7E3",
            INIT_RAM_0D => X"F6793C9E4F27B3D9DDF6793DBE4D5667C1E0E8EC3A5AAE9F93D9DDEEA753AA55B2D98CB6",
            INIT_RAM_0E => X"0A070502C26070180C06070180C06030180C06030391A8D26C860C06070A8BDAE66FB5E4",
            INIT_RAM_0F => X"0DA6BB1D8D4F6FC7E3F1F7226B66E359ACB46AC57C7E3EB67335E7F3DB8FC7633198CC4C",
            INIT_RAM_10 => X"EEE54261C0E0703865000000000000000000000000000000000000000000000097554812",
            INIT_RAM_11 => X"4A03018549E7B7D9BBF67B3D9ECF274FA7D3E9F53A9D4EA7B7A7A0F0783C1D1F06C325D4",
            INIT_RAM_12 => X"EE79E7C763B19858140A0D4501416130480C0E030180C06070180C06030189BE8EC234DA",
            INIT_RAM_13 => X"00000001900556681209367B1D8E974BC7E3F1F8F34B64E3198CB65B673C7E3EE75B43A1",
            INIT_RAM_14 => X"D0F83C1E0F0783C1516DE9558140A0502814000000000000000000000000000000000000",
            INIT_RAM_15 => X"06030381C5DF47C1D1CCD65281C4DD4FA7D3E9F9337AAEA6AB41E0F0783C1E0D872755D4",
            INIT_RAM_16 => X"6AF73C7E3E8E87ABB0CE3723B5E5F13038351AA74B49C16050461C2D88C480C0E091361C",
            INIT_RAM_17 => X"00000000000000000000000000014473381A0DB67A1D8C978FC7E3F1F7339155B3556CB6",
            INIT_RAM_18 => X"F0783C1E0F0747A3D1C9783C1E0F0783C1E0D096ABC1B0A0502814000000000000000000",
            INIT_RAM_19 => X"2E18CB20C1D151B4BB2A031769B2A2EF33E0F078332DA2A667A3D1E8F474192F06AB55E0",
            INIT_RAM_1A => X"F1F8E2B155B2D96CD5CE78FC7D2F078343D56E0494A6526130CA6532AD93A5A52850985A",
            INIT_RAM_1B => X"00000000000000000000000000000000000000000000000457AA120D84BB1D8E874BC7E3",
            INIT_RAM_1C => X"F0783C1E0F078353E0F07834150CCE8793D1D0687A3D1F074743D1E8D48B69D0A0502814",
            INIT_RAM_1D => X"52B596C9C5B194385A14000A0212A885291A8CA6D2959ACD6A35C9F0783A3E08D46BC1E0",
            INIT_RAM_1E => X"0904A33D0E86A393E3F1F8EAAD55B2D96D55F1F8FA5D1F0687AB1D092756CD6528706AB6",
            INIT_RAM_1F => X"D0F81B4140A05028140000000000000000000000000000000000000000000000CACFAC1A",
            INIT_RAM_20 => X"F0783C1E0E8D67C1E0E8F83C1E0F0783A3D1F0783A2D0001613120CCD6621A1E8F834322",
            INIT_RAM_21 => X"B7171CAB46317138D65B275AAB663318CA5B1400000001098C505AAD666B35AD0747C1E0",
            INIT_RAM_22 => X"0000000001096FAC5B09048B5A0D46ABB9E3F1F8FB8D552995B9E3F1F4BC1E0D0F54B45C",
            INIT_RAM_23 => X"0026232A988727C15159D47A25C0A0502814000000000000000000000000000000000000",
            INIT_RAM_24 => X"002633310E4F47C1E0F0783C1E0F0783C1E0F0783C1D1F0747C1E0A8EC3A3D1880000000",
            INIT_RAM_25 => X"E9783C1A2EAB7149260CB6C009B4E268005A5B2D966B65B358B6CE0C8000000000005000",
            INIT_RAM_26 => X"0000000000000000000000000001084BCF9C09048245A8CB69B8DCA6471685C2E473C7DC",
            INIT_RAM_27 => X"D8162A1C9CCC64B00000000005850A6333E0912CEA3190A0502814000000000000000000",
            INIT_RAM_28 => X"6E0640000000000000000013059906C2B3E0F0783C1D1F0747C1E0F0783C1E0F074793E0",
            INIT_RAM_29 => X"09850B8DCCDF8FA5A1F078345B42C00000191408400002CA90000059B9400E55B16DB800",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000190016D67D64D848361B2D168B614",
            INIT_RAM_2B => X"F0783C1E0F072531A1E8C8000004C381B25800000000000164B199E896D39522E050281B",
            INIT_RAM_2C => X"0037042196B270B25A00000000000000000000000005800724B1B0F0783C1E0F0783C1E0",
            INIT_RAM_2D => X"DF371345A0D068B81C0E050285C5A2CDB522A8F6E3800000000000000000000001643200",
            INIT_RAM_2E => X"A8C40329B6D050281400000000000000000000000000000000000000000000014000251C",
            INIT_RAM_2F => X"E8F83C1E0F0783C1E0F0783A3E0F07813098CCF45A000000000000000000000000000000",
            INIT_RAM_30 => X"000000000000000000000A0B2002CC9832000000000000000000000000000000034130A9",
            INIT_RAM_31 => X"0000000000000042124D5571D9ECF63AAB558AD5568B45A271CB55DA2680000000000000",
            INIT_RAM_32 => X"0000000000000000002C56400000C9702814000000000000000000000000000000000000",
            INIT_RAM_33 => X"000000000000013000ACF83C1E0F0783C1E0E8F83C1E0F078240002C4833320000000000",
            INIT_RAM_34 => X"00000000000000000000000000000000000000000000000001B600000000000000000000",
            INIT_RAM_35 => X"00000000000000000000000000000000001200064325A2D2CD66DC8E472391D8E44DB459",
            INIT_RAM_36 => X"0000000D98CA44000000000000000000000000160000000000245C000000000000000000",
            INIT_RAM_37 => X"00000000000000000000000000000000B0004C782B3D1E8F83C1E0E4F83C1D1F07839258",
            INIT_RAM_38 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_39 => X"000000000000000000000000000000000000000000000000000021001680000000000000",
            INIT_RAM_3A => X"D0727C1A0D0F83C120000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3B => X"00000000000000000000000000000000000000000000000000000014725C1D290783C1D1",
            INIT_RAM_3C => X"140000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"00441C1592C667A399D0C83C1E090687C1D12C0000000000000000000000000000000000",
            INIT_RAM_3F => X"000000000000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => promx9_inst_17_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_17,
            RESET => reset,
            AD => promx9_inst_17_AD_i
        );

    promx9_inst_18: pROMX9
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 18,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"CCA2A2144E4A27A244E4A2530C4CCA2BC183ACA2C0000000000000000000000000000000",
            INIT_RAM_05 => X"00000000000000000000000000000000000000000B0C38CB2D30C44C31130C4E4A25C0C2",
            INIT_RAM_06 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_09 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0A => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0B => X"F060E2144000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0C => X"0000000006CB2C00002C30C00007030B328A2C30E32CB4C3134285F060F328A4C313328A",
            INIT_RAM_0D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0E => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_0F => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_10 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_12 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_13 => X"8CB2CB0C328430B0C3CCA2B428590624B0C390627928954A180000000000000000000000",
            INIT_RAM_14 => X"00000000000000000000000000000000000000000000000000B0C3145280000000024189",
            INIT_RAM_15 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_16 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_18 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_19 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1A => X"00001C0C2AD32D30C4000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1B => X"00000000000000000000000000000000000054A19B2CB0000000002C30E2144CCA2A4189",
            INIT_RAM_1C => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1D => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1E => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_1F => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_20 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_21 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_22 => X"00000B0C32C30C00000000000002C30DB2CB8CB2C514A2C30DB2CB145280000000000000",
            INIT_RAM_23 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"000000000145280000000000000145280000000000000000000000000000000000000000",
            INIT_RAM_29 => X"00000B0C30000000002C30C0000145280000000000000145280000000000000145280000",
            INIT_RAM_2A => X"0000000001452800000000000001452800000000000001452800000CB14000000000514A",
            INIT_RAM_2B => X"000000000145280000000000000145280000000000000145280000000000000145280000",
            INIT_RAM_2C => X"000000000145280000000000000145280000000000000145280000000000000145280000",
            INIT_RAM_2D => X"000000000145280000000000000145280000000000000145280000000000000145280000",
            INIT_RAM_2E => X"000000000145280000000000000145280000000000000145280000000000000145280000",
            INIT_RAM_2F => X"000000000145280000000000000145280000000000000145280000000000000145280000"
        )
        port map (
            DO => promx9_inst_18_DO_o,
            CLK => clk,
            OCE => oce,
            CE => lut_f_19,
            RESET => reset,
            AD => promx9_inst_18_AD_i
        );

    dff_inst_0: DFFE
        port map (
            Q => dff_q_0,
            D => ad(14),
            CLK => clk,
            CE => ce
        );

    dff_inst_1: DFFE
        port map (
            Q => dff_q_1,
            D => ad(13),
            CLK => clk,
            CE => ce
        );

    dff_inst_2: DFFE
        port map (
            Q => dff_q_2,
            D => ad(12),
            CLK => clk,
            CE => ce
        );

    dff_inst_3: DFFE
        port map (
            Q => dff_q_3,
            D => ad(11),
            CLK => clk,
            CE => ce
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => promx9_inst_0_dout(0),
            I1 => promx9_inst_1_dout(0),
            S0 => dff_q_3
        );

    mux_inst_11: MUX2
        port map (
            O => mux_o_11,
            I0 => promx9_inst_2_dout(0),
            I1 => promx9_inst_3_dout(0),
            S0 => dff_q_3
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => promx9_inst_4_dout(0),
            I1 => promx9_inst_5_dout(0),
            S0 => dff_q_3
        );

    mux_inst_13: MUX2
        port map (
            O => mux_o_13,
            I0 => promx9_inst_6_dout(0),
            I1 => promx9_inst_7_dout(0),
            S0 => dff_q_3
        );

    mux_inst_14: MUX2
        port map (
            O => mux_o_14,
            I0 => promx9_inst_16_dout(0),
            I1 => promx9_inst_18_dout(0),
            S0 => dff_q_3
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => mux_o_10,
            I1 => mux_o_11,
            S0 => dff_q_2
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => mux_o_12,
            I1 => mux_o_13,
            S0 => dff_q_2
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => mux_o_15,
            I1 => mux_o_16,
            S0 => dff_q_1
        );

    mux_inst_20: MUX2
        port map (
            O => dout(0),
            I0 => mux_o_18,
            I1 => mux_o_14,
            S0 => dff_q_0
        );

    mux_inst_31: MUX2
        port map (
            O => mux_o_31,
            I0 => promx9_inst_0_dout(1),
            I1 => promx9_inst_1_dout(1),
            S0 => dff_q_3
        );

    mux_inst_32: MUX2
        port map (
            O => mux_o_32,
            I0 => promx9_inst_2_dout(1),
            I1 => promx9_inst_3_dout(1),
            S0 => dff_q_3
        );

    mux_inst_33: MUX2
        port map (
            O => mux_o_33,
            I0 => promx9_inst_4_dout(1),
            I1 => promx9_inst_5_dout(1),
            S0 => dff_q_3
        );

    mux_inst_34: MUX2
        port map (
            O => mux_o_34,
            I0 => promx9_inst_6_dout(1),
            I1 => promx9_inst_7_dout(1),
            S0 => dff_q_3
        );

    mux_inst_35: MUX2
        port map (
            O => mux_o_35,
            I0 => promx9_inst_16_dout(1),
            I1 => promx9_inst_18_dout(1),
            S0 => dff_q_3
        );

    mux_inst_36: MUX2
        port map (
            O => mux_o_36,
            I0 => mux_o_31,
            I1 => mux_o_32,
            S0 => dff_q_2
        );

    mux_inst_37: MUX2
        port map (
            O => mux_o_37,
            I0 => mux_o_33,
            I1 => mux_o_34,
            S0 => dff_q_2
        );

    mux_inst_39: MUX2
        port map (
            O => mux_o_39,
            I0 => mux_o_36,
            I1 => mux_o_37,
            S0 => dff_q_1
        );

    mux_inst_41: MUX2
        port map (
            O => dout(1),
            I0 => mux_o_39,
            I1 => mux_o_35,
            S0 => dff_q_0
        );

    mux_inst_52: MUX2
        port map (
            O => mux_o_52,
            I0 => promx9_inst_0_dout(2),
            I1 => promx9_inst_1_dout(2),
            S0 => dff_q_3
        );

    mux_inst_53: MUX2
        port map (
            O => mux_o_53,
            I0 => promx9_inst_2_dout(2),
            I1 => promx9_inst_3_dout(2),
            S0 => dff_q_3
        );

    mux_inst_54: MUX2
        port map (
            O => mux_o_54,
            I0 => promx9_inst_4_dout(2),
            I1 => promx9_inst_5_dout(2),
            S0 => dff_q_3
        );

    mux_inst_55: MUX2
        port map (
            O => mux_o_55,
            I0 => promx9_inst_6_dout(2),
            I1 => promx9_inst_7_dout(2),
            S0 => dff_q_3
        );

    mux_inst_56: MUX2
        port map (
            O => mux_o_56,
            I0 => promx9_inst_16_dout(2),
            I1 => promx9_inst_18_dout(2),
            S0 => dff_q_3
        );

    mux_inst_57: MUX2
        port map (
            O => mux_o_57,
            I0 => mux_o_52,
            I1 => mux_o_53,
            S0 => dff_q_2
        );

    mux_inst_58: MUX2
        port map (
            O => mux_o_58,
            I0 => mux_o_54,
            I1 => mux_o_55,
            S0 => dff_q_2
        );

    mux_inst_60: MUX2
        port map (
            O => mux_o_60,
            I0 => mux_o_57,
            I1 => mux_o_58,
            S0 => dff_q_1
        );

    mux_inst_62: MUX2
        port map (
            O => dout(2),
            I0 => mux_o_60,
            I1 => mux_o_56,
            S0 => dff_q_0
        );

    mux_inst_73: MUX2
        port map (
            O => mux_o_73,
            I0 => promx9_inst_0_dout(3),
            I1 => promx9_inst_1_dout(3),
            S0 => dff_q_3
        );

    mux_inst_74: MUX2
        port map (
            O => mux_o_74,
            I0 => promx9_inst_2_dout(3),
            I1 => promx9_inst_3_dout(3),
            S0 => dff_q_3
        );

    mux_inst_75: MUX2
        port map (
            O => mux_o_75,
            I0 => promx9_inst_4_dout(3),
            I1 => promx9_inst_5_dout(3),
            S0 => dff_q_3
        );

    mux_inst_76: MUX2
        port map (
            O => mux_o_76,
            I0 => promx9_inst_6_dout(3),
            I1 => promx9_inst_7_dout(3),
            S0 => dff_q_3
        );

    mux_inst_77: MUX2
        port map (
            O => mux_o_77,
            I0 => promx9_inst_16_dout(3),
            I1 => promx9_inst_18_dout(3),
            S0 => dff_q_3
        );

    mux_inst_78: MUX2
        port map (
            O => mux_o_78,
            I0 => mux_o_73,
            I1 => mux_o_74,
            S0 => dff_q_2
        );

    mux_inst_79: MUX2
        port map (
            O => mux_o_79,
            I0 => mux_o_75,
            I1 => mux_o_76,
            S0 => dff_q_2
        );

    mux_inst_81: MUX2
        port map (
            O => mux_o_81,
            I0 => mux_o_78,
            I1 => mux_o_79,
            S0 => dff_q_1
        );

    mux_inst_83: MUX2
        port map (
            O => dout(3),
            I0 => mux_o_81,
            I1 => mux_o_77,
            S0 => dff_q_0
        );

    mux_inst_94: MUX2
        port map (
            O => mux_o_94,
            I0 => promx9_inst_0_dout(4),
            I1 => promx9_inst_1_dout(4),
            S0 => dff_q_3
        );

    mux_inst_95: MUX2
        port map (
            O => mux_o_95,
            I0 => promx9_inst_2_dout(4),
            I1 => promx9_inst_3_dout(4),
            S0 => dff_q_3
        );

    mux_inst_96: MUX2
        port map (
            O => mux_o_96,
            I0 => promx9_inst_4_dout(4),
            I1 => promx9_inst_5_dout(4),
            S0 => dff_q_3
        );

    mux_inst_97: MUX2
        port map (
            O => mux_o_97,
            I0 => promx9_inst_6_dout(4),
            I1 => promx9_inst_7_dout(4),
            S0 => dff_q_3
        );

    mux_inst_98: MUX2
        port map (
            O => mux_o_98,
            I0 => promx9_inst_16_dout(4),
            I1 => promx9_inst_18_dout(4),
            S0 => dff_q_3
        );

    mux_inst_99: MUX2
        port map (
            O => mux_o_99,
            I0 => mux_o_94,
            I1 => mux_o_95,
            S0 => dff_q_2
        );

    mux_inst_100: MUX2
        port map (
            O => mux_o_100,
            I0 => mux_o_96,
            I1 => mux_o_97,
            S0 => dff_q_2
        );

    mux_inst_102: MUX2
        port map (
            O => mux_o_102,
            I0 => mux_o_99,
            I1 => mux_o_100,
            S0 => dff_q_1
        );

    mux_inst_104: MUX2
        port map (
            O => dout(4),
            I0 => mux_o_102,
            I1 => mux_o_98,
            S0 => dff_q_0
        );

    mux_inst_115: MUX2
        port map (
            O => mux_o_115,
            I0 => promx9_inst_0_dout(5),
            I1 => promx9_inst_1_dout(5),
            S0 => dff_q_3
        );

    mux_inst_116: MUX2
        port map (
            O => mux_o_116,
            I0 => promx9_inst_2_dout(5),
            I1 => promx9_inst_3_dout(5),
            S0 => dff_q_3
        );

    mux_inst_117: MUX2
        port map (
            O => mux_o_117,
            I0 => promx9_inst_4_dout(5),
            I1 => promx9_inst_5_dout(5),
            S0 => dff_q_3
        );

    mux_inst_118: MUX2
        port map (
            O => mux_o_118,
            I0 => promx9_inst_6_dout(5),
            I1 => promx9_inst_7_dout(5),
            S0 => dff_q_3
        );

    mux_inst_119: MUX2
        port map (
            O => mux_o_119,
            I0 => promx9_inst_16_dout(5),
            I1 => promx9_inst_18_dout(5),
            S0 => dff_q_3
        );

    mux_inst_120: MUX2
        port map (
            O => mux_o_120,
            I0 => mux_o_115,
            I1 => mux_o_116,
            S0 => dff_q_2
        );

    mux_inst_121: MUX2
        port map (
            O => mux_o_121,
            I0 => mux_o_117,
            I1 => mux_o_118,
            S0 => dff_q_2
        );

    mux_inst_123: MUX2
        port map (
            O => mux_o_123,
            I0 => mux_o_120,
            I1 => mux_o_121,
            S0 => dff_q_1
        );

    mux_inst_125: MUX2
        port map (
            O => dout(5),
            I0 => mux_o_123,
            I1 => mux_o_119,
            S0 => dff_q_0
        );

    mux_inst_136: MUX2
        port map (
            O => mux_o_136,
            I0 => promx9_inst_0_dout(6),
            I1 => promx9_inst_1_dout(6),
            S0 => dff_q_3
        );

    mux_inst_137: MUX2
        port map (
            O => mux_o_137,
            I0 => promx9_inst_2_dout(6),
            I1 => promx9_inst_3_dout(6),
            S0 => dff_q_3
        );

    mux_inst_138: MUX2
        port map (
            O => mux_o_138,
            I0 => promx9_inst_4_dout(6),
            I1 => promx9_inst_5_dout(6),
            S0 => dff_q_3
        );

    mux_inst_139: MUX2
        port map (
            O => mux_o_139,
            I0 => promx9_inst_6_dout(6),
            I1 => promx9_inst_7_dout(6),
            S0 => dff_q_3
        );

    mux_inst_140: MUX2
        port map (
            O => mux_o_140,
            I0 => promx9_inst_16_dout(6),
            I1 => promx9_inst_18_dout(6),
            S0 => dff_q_3
        );

    mux_inst_141: MUX2
        port map (
            O => mux_o_141,
            I0 => mux_o_136,
            I1 => mux_o_137,
            S0 => dff_q_2
        );

    mux_inst_142: MUX2
        port map (
            O => mux_o_142,
            I0 => mux_o_138,
            I1 => mux_o_139,
            S0 => dff_q_2
        );

    mux_inst_144: MUX2
        port map (
            O => mux_o_144,
            I0 => mux_o_141,
            I1 => mux_o_142,
            S0 => dff_q_1
        );

    mux_inst_146: MUX2
        port map (
            O => dout(6),
            I0 => mux_o_144,
            I1 => mux_o_140,
            S0 => dff_q_0
        );

    mux_inst_157: MUX2
        port map (
            O => mux_o_157,
            I0 => promx9_inst_0_dout(7),
            I1 => promx9_inst_1_dout(7),
            S0 => dff_q_3
        );

    mux_inst_158: MUX2
        port map (
            O => mux_o_158,
            I0 => promx9_inst_2_dout(7),
            I1 => promx9_inst_3_dout(7),
            S0 => dff_q_3
        );

    mux_inst_159: MUX2
        port map (
            O => mux_o_159,
            I0 => promx9_inst_4_dout(7),
            I1 => promx9_inst_5_dout(7),
            S0 => dff_q_3
        );

    mux_inst_160: MUX2
        port map (
            O => mux_o_160,
            I0 => promx9_inst_6_dout(7),
            I1 => promx9_inst_7_dout(7),
            S0 => dff_q_3
        );

    mux_inst_161: MUX2
        port map (
            O => mux_o_161,
            I0 => promx9_inst_16_dout(7),
            I1 => promx9_inst_18_dout(7),
            S0 => dff_q_3
        );

    mux_inst_162: MUX2
        port map (
            O => mux_o_162,
            I0 => mux_o_157,
            I1 => mux_o_158,
            S0 => dff_q_2
        );

    mux_inst_163: MUX2
        port map (
            O => mux_o_163,
            I0 => mux_o_159,
            I1 => mux_o_160,
            S0 => dff_q_2
        );

    mux_inst_165: MUX2
        port map (
            O => mux_o_165,
            I0 => mux_o_162,
            I1 => mux_o_163,
            S0 => dff_q_1
        );

    mux_inst_167: MUX2
        port map (
            O => dout(7),
            I0 => mux_o_165,
            I1 => mux_o_161,
            S0 => dff_q_0
        );

    mux_inst_178: MUX2
        port map (
            O => mux_o_178,
            I0 => promx9_inst_0_dout(8),
            I1 => promx9_inst_1_dout(8),
            S0 => dff_q_3
        );

    mux_inst_179: MUX2
        port map (
            O => mux_o_179,
            I0 => promx9_inst_2_dout(8),
            I1 => promx9_inst_3_dout(8),
            S0 => dff_q_3
        );

    mux_inst_180: MUX2
        port map (
            O => mux_o_180,
            I0 => promx9_inst_4_dout(8),
            I1 => promx9_inst_5_dout(8),
            S0 => dff_q_3
        );

    mux_inst_181: MUX2
        port map (
            O => mux_o_181,
            I0 => promx9_inst_6_dout(8),
            I1 => promx9_inst_7_dout(8),
            S0 => dff_q_3
        );

    mux_inst_182: MUX2
        port map (
            O => mux_o_182,
            I0 => promx9_inst_16_dout(8),
            I1 => promx9_inst_18_dout(8),
            S0 => dff_q_3
        );

    mux_inst_183: MUX2
        port map (
            O => mux_o_183,
            I0 => mux_o_178,
            I1 => mux_o_179,
            S0 => dff_q_2
        );

    mux_inst_184: MUX2
        port map (
            O => mux_o_184,
            I0 => mux_o_180,
            I1 => mux_o_181,
            S0 => dff_q_2
        );

    mux_inst_186: MUX2
        port map (
            O => mux_o_186,
            I0 => mux_o_183,
            I1 => mux_o_184,
            S0 => dff_q_1
        );

    mux_inst_188: MUX2
        port map (
            O => dout(8),
            I0 => mux_o_186,
            I1 => mux_o_182,
            S0 => dff_q_0
        );

    mux_inst_199: MUX2
        port map (
            O => mux_o_199,
            I0 => promx9_inst_8_dout(9),
            I1 => promx9_inst_9_dout(9),
            S0 => dff_q_3
        );

    mux_inst_200: MUX2
        port map (
            O => mux_o_200,
            I0 => promx9_inst_10_dout(9),
            I1 => promx9_inst_11_dout(9),
            S0 => dff_q_3
        );

    mux_inst_201: MUX2
        port map (
            O => mux_o_201,
            I0 => promx9_inst_12_dout(9),
            I1 => promx9_inst_13_dout(9),
            S0 => dff_q_3
        );

    mux_inst_202: MUX2
        port map (
            O => mux_o_202,
            I0 => promx9_inst_14_dout(9),
            I1 => promx9_inst_15_dout(9),
            S0 => dff_q_3
        );

    mux_inst_203: MUX2
        port map (
            O => mux_o_203,
            I0 => promx9_inst_17_dout(9),
            I1 => promx9_inst_18_dout(9),
            S0 => dff_q_3
        );

    mux_inst_204: MUX2
        port map (
            O => mux_o_204,
            I0 => mux_o_199,
            I1 => mux_o_200,
            S0 => dff_q_2
        );

    mux_inst_205: MUX2
        port map (
            O => mux_o_205,
            I0 => mux_o_201,
            I1 => mux_o_202,
            S0 => dff_q_2
        );

    mux_inst_207: MUX2
        port map (
            O => mux_o_207,
            I0 => mux_o_204,
            I1 => mux_o_205,
            S0 => dff_q_1
        );

    mux_inst_209: MUX2
        port map (
            O => dout(9),
            I0 => mux_o_207,
            I1 => mux_o_203,
            S0 => dff_q_0
        );

    mux_inst_220: MUX2
        port map (
            O => mux_o_220,
            I0 => promx9_inst_8_dout(10),
            I1 => promx9_inst_9_dout(10),
            S0 => dff_q_3
        );

    mux_inst_221: MUX2
        port map (
            O => mux_o_221,
            I0 => promx9_inst_10_dout(10),
            I1 => promx9_inst_11_dout(10),
            S0 => dff_q_3
        );

    mux_inst_222: MUX2
        port map (
            O => mux_o_222,
            I0 => promx9_inst_12_dout(10),
            I1 => promx9_inst_13_dout(10),
            S0 => dff_q_3
        );

    mux_inst_223: MUX2
        port map (
            O => mux_o_223,
            I0 => promx9_inst_14_dout(10),
            I1 => promx9_inst_15_dout(10),
            S0 => dff_q_3
        );

    mux_inst_224: MUX2
        port map (
            O => mux_o_224,
            I0 => promx9_inst_17_dout(10),
            I1 => promx9_inst_18_dout(10),
            S0 => dff_q_3
        );

    mux_inst_225: MUX2
        port map (
            O => mux_o_225,
            I0 => mux_o_220,
            I1 => mux_o_221,
            S0 => dff_q_2
        );

    mux_inst_226: MUX2
        port map (
            O => mux_o_226,
            I0 => mux_o_222,
            I1 => mux_o_223,
            S0 => dff_q_2
        );

    mux_inst_228: MUX2
        port map (
            O => mux_o_228,
            I0 => mux_o_225,
            I1 => mux_o_226,
            S0 => dff_q_1
        );

    mux_inst_230: MUX2
        port map (
            O => dout(10),
            I0 => mux_o_228,
            I1 => mux_o_224,
            S0 => dff_q_0
        );

    mux_inst_241: MUX2
        port map (
            O => mux_o_241,
            I0 => promx9_inst_8_dout(11),
            I1 => promx9_inst_9_dout(11),
            S0 => dff_q_3
        );

    mux_inst_242: MUX2
        port map (
            O => mux_o_242,
            I0 => promx9_inst_10_dout(11),
            I1 => promx9_inst_11_dout(11),
            S0 => dff_q_3
        );

    mux_inst_243: MUX2
        port map (
            O => mux_o_243,
            I0 => promx9_inst_12_dout(11),
            I1 => promx9_inst_13_dout(11),
            S0 => dff_q_3
        );

    mux_inst_244: MUX2
        port map (
            O => mux_o_244,
            I0 => promx9_inst_14_dout(11),
            I1 => promx9_inst_15_dout(11),
            S0 => dff_q_3
        );

    mux_inst_245: MUX2
        port map (
            O => mux_o_245,
            I0 => promx9_inst_17_dout(11),
            I1 => promx9_inst_18_dout(11),
            S0 => dff_q_3
        );

    mux_inst_246: MUX2
        port map (
            O => mux_o_246,
            I0 => mux_o_241,
            I1 => mux_o_242,
            S0 => dff_q_2
        );

    mux_inst_247: MUX2
        port map (
            O => mux_o_247,
            I0 => mux_o_243,
            I1 => mux_o_244,
            S0 => dff_q_2
        );

    mux_inst_249: MUX2
        port map (
            O => mux_o_249,
            I0 => mux_o_246,
            I1 => mux_o_247,
            S0 => dff_q_1
        );

    mux_inst_251: MUX2
        port map (
            O => dout(11),
            I0 => mux_o_249,
            I1 => mux_o_245,
            S0 => dff_q_0
        );

    mux_inst_262: MUX2
        port map (
            O => mux_o_262,
            I0 => promx9_inst_8_dout(12),
            I1 => promx9_inst_9_dout(12),
            S0 => dff_q_3
        );

    mux_inst_263: MUX2
        port map (
            O => mux_o_263,
            I0 => promx9_inst_10_dout(12),
            I1 => promx9_inst_11_dout(12),
            S0 => dff_q_3
        );

    mux_inst_264: MUX2
        port map (
            O => mux_o_264,
            I0 => promx9_inst_12_dout(12),
            I1 => promx9_inst_13_dout(12),
            S0 => dff_q_3
        );

    mux_inst_265: MUX2
        port map (
            O => mux_o_265,
            I0 => promx9_inst_14_dout(12),
            I1 => promx9_inst_15_dout(12),
            S0 => dff_q_3
        );

    mux_inst_266: MUX2
        port map (
            O => mux_o_266,
            I0 => promx9_inst_17_dout(12),
            I1 => promx9_inst_18_dout(12),
            S0 => dff_q_3
        );

    mux_inst_267: MUX2
        port map (
            O => mux_o_267,
            I0 => mux_o_262,
            I1 => mux_o_263,
            S0 => dff_q_2
        );

    mux_inst_268: MUX2
        port map (
            O => mux_o_268,
            I0 => mux_o_264,
            I1 => mux_o_265,
            S0 => dff_q_2
        );

    mux_inst_270: MUX2
        port map (
            O => mux_o_270,
            I0 => mux_o_267,
            I1 => mux_o_268,
            S0 => dff_q_1
        );

    mux_inst_272: MUX2
        port map (
            O => dout(12),
            I0 => mux_o_270,
            I1 => mux_o_266,
            S0 => dff_q_0
        );

    mux_inst_283: MUX2
        port map (
            O => mux_o_283,
            I0 => promx9_inst_8_dout(13),
            I1 => promx9_inst_9_dout(13),
            S0 => dff_q_3
        );

    mux_inst_284: MUX2
        port map (
            O => mux_o_284,
            I0 => promx9_inst_10_dout(13),
            I1 => promx9_inst_11_dout(13),
            S0 => dff_q_3
        );

    mux_inst_285: MUX2
        port map (
            O => mux_o_285,
            I0 => promx9_inst_12_dout(13),
            I1 => promx9_inst_13_dout(13),
            S0 => dff_q_3
        );

    mux_inst_286: MUX2
        port map (
            O => mux_o_286,
            I0 => promx9_inst_14_dout(13),
            I1 => promx9_inst_15_dout(13),
            S0 => dff_q_3
        );

    mux_inst_287: MUX2
        port map (
            O => mux_o_287,
            I0 => promx9_inst_17_dout(13),
            I1 => promx9_inst_18_dout(13),
            S0 => dff_q_3
        );

    mux_inst_288: MUX2
        port map (
            O => mux_o_288,
            I0 => mux_o_283,
            I1 => mux_o_284,
            S0 => dff_q_2
        );

    mux_inst_289: MUX2
        port map (
            O => mux_o_289,
            I0 => mux_o_285,
            I1 => mux_o_286,
            S0 => dff_q_2
        );

    mux_inst_291: MUX2
        port map (
            O => mux_o_291,
            I0 => mux_o_288,
            I1 => mux_o_289,
            S0 => dff_q_1
        );

    mux_inst_293: MUX2
        port map (
            O => dout(13),
            I0 => mux_o_291,
            I1 => mux_o_287,
            S0 => dff_q_0
        );

    mux_inst_304: MUX2
        port map (
            O => mux_o_304,
            I0 => promx9_inst_8_dout(14),
            I1 => promx9_inst_9_dout(14),
            S0 => dff_q_3
        );

    mux_inst_305: MUX2
        port map (
            O => mux_o_305,
            I0 => promx9_inst_10_dout(14),
            I1 => promx9_inst_11_dout(14),
            S0 => dff_q_3
        );

    mux_inst_306: MUX2
        port map (
            O => mux_o_306,
            I0 => promx9_inst_12_dout(14),
            I1 => promx9_inst_13_dout(14),
            S0 => dff_q_3
        );

    mux_inst_307: MUX2
        port map (
            O => mux_o_307,
            I0 => promx9_inst_14_dout(14),
            I1 => promx9_inst_15_dout(14),
            S0 => dff_q_3
        );

    mux_inst_308: MUX2
        port map (
            O => mux_o_308,
            I0 => promx9_inst_17_dout(14),
            I1 => promx9_inst_18_dout(14),
            S0 => dff_q_3
        );

    mux_inst_309: MUX2
        port map (
            O => mux_o_309,
            I0 => mux_o_304,
            I1 => mux_o_305,
            S0 => dff_q_2
        );

    mux_inst_310: MUX2
        port map (
            O => mux_o_310,
            I0 => mux_o_306,
            I1 => mux_o_307,
            S0 => dff_q_2
        );

    mux_inst_312: MUX2
        port map (
            O => mux_o_312,
            I0 => mux_o_309,
            I1 => mux_o_310,
            S0 => dff_q_1
        );

    mux_inst_314: MUX2
        port map (
            O => dout(14),
            I0 => mux_o_312,
            I1 => mux_o_308,
            S0 => dff_q_0
        );

    mux_inst_325: MUX2
        port map (
            O => mux_o_325,
            I0 => promx9_inst_8_dout(15),
            I1 => promx9_inst_9_dout(15),
            S0 => dff_q_3
        );

    mux_inst_326: MUX2
        port map (
            O => mux_o_326,
            I0 => promx9_inst_10_dout(15),
            I1 => promx9_inst_11_dout(15),
            S0 => dff_q_3
        );

    mux_inst_327: MUX2
        port map (
            O => mux_o_327,
            I0 => promx9_inst_12_dout(15),
            I1 => promx9_inst_13_dout(15),
            S0 => dff_q_3
        );

    mux_inst_328: MUX2
        port map (
            O => mux_o_328,
            I0 => promx9_inst_14_dout(15),
            I1 => promx9_inst_15_dout(15),
            S0 => dff_q_3
        );

    mux_inst_329: MUX2
        port map (
            O => mux_o_329,
            I0 => promx9_inst_17_dout(15),
            I1 => promx9_inst_18_dout(15),
            S0 => dff_q_3
        );

    mux_inst_330: MUX2
        port map (
            O => mux_o_330,
            I0 => mux_o_325,
            I1 => mux_o_326,
            S0 => dff_q_2
        );

    mux_inst_331: MUX2
        port map (
            O => mux_o_331,
            I0 => mux_o_327,
            I1 => mux_o_328,
            S0 => dff_q_2
        );

    mux_inst_333: MUX2
        port map (
            O => mux_o_333,
            I0 => mux_o_330,
            I1 => mux_o_331,
            S0 => dff_q_1
        );

    mux_inst_335: MUX2
        port map (
            O => dout(15),
            I0 => mux_o_333,
            I1 => mux_o_329,
            S0 => dff_q_0
        );

    mux_inst_346: MUX2
        port map (
            O => mux_o_346,
            I0 => promx9_inst_8_dout(16),
            I1 => promx9_inst_9_dout(16),
            S0 => dff_q_3
        );

    mux_inst_347: MUX2
        port map (
            O => mux_o_347,
            I0 => promx9_inst_10_dout(16),
            I1 => promx9_inst_11_dout(16),
            S0 => dff_q_3
        );

    mux_inst_348: MUX2
        port map (
            O => mux_o_348,
            I0 => promx9_inst_12_dout(16),
            I1 => promx9_inst_13_dout(16),
            S0 => dff_q_3
        );

    mux_inst_349: MUX2
        port map (
            O => mux_o_349,
            I0 => promx9_inst_14_dout(16),
            I1 => promx9_inst_15_dout(16),
            S0 => dff_q_3
        );

    mux_inst_350: MUX2
        port map (
            O => mux_o_350,
            I0 => promx9_inst_17_dout(16),
            I1 => promx9_inst_18_dout(16),
            S0 => dff_q_3
        );

    mux_inst_351: MUX2
        port map (
            O => mux_o_351,
            I0 => mux_o_346,
            I1 => mux_o_347,
            S0 => dff_q_2
        );

    mux_inst_352: MUX2
        port map (
            O => mux_o_352,
            I0 => mux_o_348,
            I1 => mux_o_349,
            S0 => dff_q_2
        );

    mux_inst_354: MUX2
        port map (
            O => mux_o_354,
            I0 => mux_o_351,
            I1 => mux_o_352,
            S0 => dff_q_1
        );

    mux_inst_356: MUX2
        port map (
            O => dout(16),
            I0 => mux_o_354,
            I1 => mux_o_350,
            S0 => dff_q_0
        );

    mux_inst_367: MUX2
        port map (
            O => mux_o_367,
            I0 => promx9_inst_8_dout(17),
            I1 => promx9_inst_9_dout(17),
            S0 => dff_q_3
        );

    mux_inst_368: MUX2
        port map (
            O => mux_o_368,
            I0 => promx9_inst_10_dout(17),
            I1 => promx9_inst_11_dout(17),
            S0 => dff_q_3
        );

    mux_inst_369: MUX2
        port map (
            O => mux_o_369,
            I0 => promx9_inst_12_dout(17),
            I1 => promx9_inst_13_dout(17),
            S0 => dff_q_3
        );

    mux_inst_370: MUX2
        port map (
            O => mux_o_370,
            I0 => promx9_inst_14_dout(17),
            I1 => promx9_inst_15_dout(17),
            S0 => dff_q_3
        );

    mux_inst_371: MUX2
        port map (
            O => mux_o_371,
            I0 => promx9_inst_17_dout(17),
            I1 => promx9_inst_18_dout(17),
            S0 => dff_q_3
        );

    mux_inst_372: MUX2
        port map (
            O => mux_o_372,
            I0 => mux_o_367,
            I1 => mux_o_368,
            S0 => dff_q_2
        );

    mux_inst_373: MUX2
        port map (
            O => mux_o_373,
            I0 => mux_o_369,
            I1 => mux_o_370,
            S0 => dff_q_2
        );

    mux_inst_375: MUX2
        port map (
            O => mux_o_375,
            I0 => mux_o_372,
            I1 => mux_o_373,
            S0 => dff_q_1
        );

    mux_inst_377: MUX2
        port map (
            O => dout(17),
            I0 => mux_o_375,
            I1 => mux_o_371,
            S0 => dff_q_0
        );

end Behavioral; --gato_colorido
